// CurrCTRL_SYS.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module CurrCTRL_SYS (
		input  wire        clk_currctrl_sys_fifo_clk,                   //           clk_currctrl_sys_fifo.clk
		input  wire        clk_currctrl_sys_ram_clk,                    //            clk_currctrl_sys_ram.clk
		input  wire        clk_pheripal_clk,                            //                    clk_pheripal.clk
		input  wire        cpu_clk_clk,                                 //                         cpu_clk.clk
		input  wire        cpu_reset_reset_n,                           //                       cpu_reset.reset_n
		input  wire [31:0] currctrl_gpio_ext_in_port,                   //               currctrl_gpio_ext.in_port
		output wire [31:0] currctrl_gpio_ext_out_port,                  //                                .out_port
		input  wire [2:0]  currctrl_gpio_s1_address,                    //                currctrl_gpio_s1.address
		input  wire        currctrl_gpio_s1_write_n,                    //                                .write_n
		input  wire [31:0] currctrl_gpio_s1_writedata,                  //                                .writedata
		input  wire        currctrl_gpio_s1_chipselect,                 //                                .chipselect
		output wire [31:0] currctrl_gpio_s1_readdata,                   //                                .readdata
		input  wire [7:0]  currctrl_register_ram_s1_address,            //        currctrl_register_ram_s1.address
		input  wire        currctrl_register_ram_s1_clken,              //                                .clken
		input  wire        currctrl_register_ram_s1_chipselect,         //                                .chipselect
		input  wire        currctrl_register_ram_s1_write,              //                                .write
		output wire [31:0] currctrl_register_ram_s1_readdata,           //                                .readdata
		input  wire [31:0] currctrl_register_ram_s1_writedata,          //                                .writedata
		input  wire [3:0]  currctrl_register_ram_s1_byteenable,         //                                .byteenable
		input  wire [7:0]  currctrl_register_ram_s2_address,            //        currctrl_register_ram_s2.address
		input  wire        currctrl_register_ram_s2_chipselect,         //                                .chipselect
		input  wire        currctrl_register_ram_s2_clken,              //                                .clken
		input  wire        currctrl_register_ram_s2_write,              //                                .write
		output wire [31:0] currctrl_register_ram_s2_readdata,           //                                .readdata
		input  wire [31:0] currctrl_register_ram_s2_writedata,          //                                .writedata
		input  wire [3:0]  currctrl_register_ram_s2_byteenable,         //                                .byteenable
		input  wire        currctrlsys_bridge_acknowledge,              //              currctrlsys_bridge.acknowledge
		input  wire        currctrlsys_bridge_irq,                      //                                .irq
		output wire [6:0]  currctrlsys_bridge_address,                  //                                .address
		output wire        currctrlsys_bridge_bus_enable,               //                                .bus_enable
		output wire [3:0]  currctrlsys_bridge_byte_enable,              //                                .byte_enable
		output wire        currctrlsys_bridge_rw,                       //                                .rw
		output wire [31:0] currctrlsys_bridge_write_data,               //                                .write_data
		input  wire [31:0] currctrlsys_bridge_read_data,                //                                .read_data
		input  wire [4:0]  currctrlsys_bridge_avalon_slave_address,     // currctrlsys_bridge_avalon_slave.address
		input  wire [3:0]  currctrlsys_bridge_avalon_slave_byteenable,  //                                .byteenable
		input  wire        currctrlsys_bridge_avalon_slave_chipselect,  //                                .chipselect
		input  wire        currctrlsys_bridge_avalon_slave_read,        //                                .read
		input  wire        currctrlsys_bridge_avalon_slave_write,       //                                .write
		input  wire [31:0] currctrlsys_bridge_avalon_slave_writedata,   //                                .writedata
		output wire [31:0] currctrlsys_bridge_avalon_slave_readdata,    //                                .readdata
		output wire        currctrlsys_bridge_avalon_slave_waitrequest, //                                .waitrequest
		output wire        currctrlsys_bridge_interrupt_irq,            //    currctrlsys_bridge_interrupt.irq
		input  wire        reset_currctrl_sys_fifo_reset_n,             //         reset_currctrl_sys_fifo.reset_n
		input  wire        reset_currctrl_sys_ram_reset_n,              //          reset_currctrl_sys_ram.reset_n
		input  wire        reset_pheripal_reset_n                       //                  reset_pheripal.reset_n
	);

	wire    rst_controller_reset_out_reset;         // rst_controller:reset_out -> [CurrCTRLSYS_Bridge:reset, CurrCTRL_GPIO:reset_n, CurrCTRL_Register_RAM:reset]
	wire    rst_controller_reset_out_reset_req;     // rst_controller:reset_req -> [CurrCTRL_Register_RAM:reset_req, rst_translator:reset_req_in]
	wire    rst_controller_001_reset_out_reset;     // rst_controller_001:reset_out -> CurrCTRL_Register_RAM:reset2
	wire    rst_controller_001_reset_out_reset_req; // rst_controller_001:reset_req -> CurrCTRL_Register_RAM:reset_req2

	CurrCTRL_SYS_CurrCTRLSYS_Bridge currctrlsys_bridge (
		.clk                (clk_pheripal_clk),                            //                clk.clk
		.reset              (rst_controller_reset_out_reset),              //              reset.reset
		.avalon_address     (currctrlsys_bridge_avalon_slave_address),     //       avalon_slave.address
		.avalon_byteenable  (currctrlsys_bridge_avalon_slave_byteenable),  //                   .byteenable
		.avalon_chipselect  (currctrlsys_bridge_avalon_slave_chipselect),  //                   .chipselect
		.avalon_read        (currctrlsys_bridge_avalon_slave_read),        //                   .read
		.avalon_write       (currctrlsys_bridge_avalon_slave_write),       //                   .write
		.avalon_writedata   (currctrlsys_bridge_avalon_slave_writedata),   //                   .writedata
		.avalon_readdata    (currctrlsys_bridge_avalon_slave_readdata),    //                   .readdata
		.avalon_waitrequest (currctrlsys_bridge_avalon_slave_waitrequest), //                   .waitrequest
		.avalon_irq         (currctrlsys_bridge_interrupt_irq),            //          interrupt.irq
		.acknowledge        (currctrlsys_bridge_acknowledge),              // external_interface.export
		.irq                (currctrlsys_bridge_irq),                      //                   .export
		.address            (currctrlsys_bridge_address),                  //                   .export
		.bus_enable         (currctrlsys_bridge_bus_enable),               //                   .export
		.byte_enable        (currctrlsys_bridge_byte_enable),              //                   .export
		.rw                 (currctrlsys_bridge_rw),                       //                   .export
		.write_data         (currctrlsys_bridge_write_data),               //                   .export
		.read_data          (currctrlsys_bridge_read_data)                 //                   .export
	);

	CurrCTRL_SYS_CurrCTRL_GPIO currctrl_gpio (
		.clk        (clk_pheripal_clk),                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset), //               reset.reset_n
		.address    (currctrl_gpio_s1_address),        //                  s1.address
		.write_n    (currctrl_gpio_s1_write_n),        //                    .write_n
		.writedata  (currctrl_gpio_s1_writedata),      //                    .writedata
		.chipselect (currctrl_gpio_s1_chipselect),     //                    .chipselect
		.readdata   (currctrl_gpio_s1_readdata),       //                    .readdata
		.in_port    (currctrl_gpio_ext_in_port),       // external_connection.export
		.out_port   (currctrl_gpio_ext_out_port)       //                    .export
	);

	CurrCTRL_SYS_CurrCTRL_Register_RAM currctrl_register_ram (
		.clk         (clk_pheripal_clk),                       //   clk1.clk
		.address     (currctrl_register_ram_s1_address),       //     s1.address
		.clken       (currctrl_register_ram_s1_clken),         //       .clken
		.chipselect  (currctrl_register_ram_s1_chipselect),    //       .chipselect
		.write       (currctrl_register_ram_s1_write),         //       .write
		.readdata    (currctrl_register_ram_s1_readdata),      //       .readdata
		.writedata   (currctrl_register_ram_s1_writedata),     //       .writedata
		.byteenable  (currctrl_register_ram_s1_byteenable),    //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.address2    (currctrl_register_ram_s2_address),       //     s2.address
		.chipselect2 (currctrl_register_ram_s2_chipselect),    //       .chipselect
		.clken2      (currctrl_register_ram_s2_clken),         //       .clken
		.write2      (currctrl_register_ram_s2_write),         //       .write
		.readdata2   (currctrl_register_ram_s2_readdata),      //       .readdata
		.writedata2  (currctrl_register_ram_s2_writedata),     //       .writedata
		.byteenable2 (currctrl_register_ram_s2_byteenable),    //       .byteenable
		.clk2        (clk_currctrl_sys_fifo_clk),              //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_pheripal_reset_n),            // reset_in0.reset
		.clk            (clk_pheripal_clk),                   //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_currctrl_sys_fifo_reset_n),       // reset_in0.reset
		.clk            (clk_currctrl_sys_fifo_clk),              //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
