
module pll_2 (
	altpll_0_locked_conduit_export,
	clk_clk,
	clk_200m_clk,
	clk_50m_clk,
	reset_reset_n);	

	output		altpll_0_locked_conduit_export;
	input		clk_clk;
	output		clk_200m_clk;
	output		clk_50m_clk;
	input		reset_reset_n;
endmodule
