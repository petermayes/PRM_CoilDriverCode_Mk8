// Mk8_InlineController_CPU_PatternGeneratorSYS_0.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module Mk8_InlineController_CPU_PatternGeneratorSYS_0 (
		input  wire        pd_clk_clk,                //          pd_clk.clk
		input  wire [3:0]  pd_debugram_s1_address,    //  pd_debugram_s1.address
		input  wire        pd_debugram_s1_clken,      //                .clken
		input  wire        pd_debugram_s1_chipselect, //                .chipselect
		input  wire        pd_debugram_s1_write,      //                .write
		output wire [31:0] pd_debugram_s1_readdata,   //                .readdata
		input  wire [31:0] pd_debugram_s1_writedata,  //                .writedata
		input  wire [3:0]  pd_debugram_s1_byteenable, //                .byteenable
		input  wire [3:0]  pd_debugram_s2_address,    //  pd_debugram_s2.address
		input  wire        pd_debugram_s2_chipselect, //                .chipselect
		input  wire        pd_debugram_s2_clken,      //                .clken
		input  wire        pd_debugram_s2_write,      //                .write
		output wire [31:0] pd_debugram_s2_readdata,   //                .readdata
		input  wire [31:0] pd_debugram_s2_writedata,  //                .writedata
		input  wire [3:0]  pd_debugram_s2_byteenable, //                .byteenable
		input  wire [31:0] pd_fifo_in_writedata,      //      pd_fifo_in.writedata
		input  wire        pd_fifo_in_write,          //                .write
		output wire        pd_fifo_in_waitrequest,    //                .waitrequest
		input  wire [2:0]  pd_fifo_in_csr_address,    //  pd_fifo_in_csr.address
		input  wire        pd_fifo_in_csr_read,       //                .read
		input  wire [31:0] pd_fifo_in_csr_writedata,  //                .writedata
		input  wire        pd_fifo_in_csr_write,      //                .write
		output wire [31:0] pd_fifo_in_csr_readdata,   //                .readdata
		output wire [31:0] pd_fifo_out_readdata,      //     pd_fifo_out.readdata
		input  wire        pd_fifo_out_read,          //                .read
		output wire        pd_fifo_out_waitrequest,   //                .waitrequest
		input  wire [2:0]  pd_fifo_out_csr_address,   // pd_fifo_out_csr.address
		input  wire        pd_fifo_out_csr_read,      //                .read
		input  wire [31:0] pd_fifo_out_csr_writedata, //                .writedata
		input  wire        pd_fifo_out_csr_write,     //                .write
		output wire [31:0] pd_fifo_out_csr_readdata,  //                .readdata
		input  wire [31:0] pd_gpio_in_port,           //         pd_gpio.in_port
		output wire [31:0] pd_gpio_out_port,          //                .out_port
		input  wire [2:0]  pd_gpio_s1_address,        //      pd_gpio_s1.address
		input  wire        pd_gpio_s1_write_n,        //                .write_n
		input  wire [31:0] pd_gpio_s1_writedata,      //                .writedata
		input  wire        pd_gpio_s1_chipselect,     //                .chipselect
		output wire [31:0] pd_gpio_s1_readdata,       //                .readdata
		input  wire        pd_reset_reset_n,          //        pd_reset.reset_n
		input  wire        pheriphal_clk_clk,         //   pheriphal_clk.clk
		input  wire        pheriphal_reset_reset_n,   // pheriphal_reset.reset_n
		output wire        reset_out_export,          //       reset_out.export
		input  wire [2:0]  reset_pd_s1_address,       //     reset_pd_s1.address
		input  wire        reset_pd_s1_write_n,       //                .write_n
		input  wire [31:0] reset_pd_s1_writedata,     //                .writedata
		input  wire        reset_pd_s1_chipselect,    //                .chipselect
		output wire [31:0] reset_pd_s1_readdata       //                .readdata
	);

	wire    rst_controller_reset_out_reset;         // rst_controller:reset_out -> [PD_DebugRAM:reset, PD_FIFO:wrreset_n, PD_GPIO:reset_n, Reset_PD:reset_n, rst_translator:in_reset]
	wire    rst_controller_reset_out_reset_req;     // rst_controller:reset_req -> [PD_DebugRAM:reset_req, rst_translator:reset_req_in]
	wire    rst_controller_001_reset_out_reset;     // rst_controller_001:reset_out -> [PD_DebugRAM:reset2, PD_FIFO:rdreset_n]
	wire    rst_controller_001_reset_out_reset_req; // rst_controller_001:reset_req -> PD_DebugRAM:reset_req2

	Mk8_InlineController_CPU_PatternGeneratorSYS_0_PD_DebugRAM pd_debugram (
		.clk         (pheriphal_clk_clk),                      //   clk1.clk
		.address     (pd_debugram_s1_address),                 //     s1.address
		.clken       (pd_debugram_s1_clken),                   //       .clken
		.chipselect  (pd_debugram_s1_chipselect),              //       .chipselect
		.write       (pd_debugram_s1_write),                   //       .write
		.readdata    (pd_debugram_s1_readdata),                //       .readdata
		.writedata   (pd_debugram_s1_writedata),               //       .writedata
		.byteenable  (pd_debugram_s1_byteenable),              //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.address2    (pd_debugram_s2_address),                 //     s2.address
		.chipselect2 (pd_debugram_s2_chipselect),              //       .chipselect
		.clken2      (pd_debugram_s2_clken),                   //       .clken
		.write2      (pd_debugram_s2_write),                   //       .write
		.readdata2   (pd_debugram_s2_readdata),                //       .readdata
		.writedata2  (pd_debugram_s2_writedata),               //       .writedata
		.byteenable2 (pd_debugram_s2_byteenable),              //       .byteenable
		.clk2        (pd_clk_clk),                             //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	Mk8_InlineController_CPU_PatternGeneratorSYS_0_PD_FIFO pd_fifo (
		.wrclock                          (pheriphal_clk_clk),                   //    clk_in.clk
		.wrreset_n                        (~rst_controller_reset_out_reset),     //  reset_in.reset_n
		.rdclock                          (pd_clk_clk),                          //   clk_out.clk
		.rdreset_n                        (~rst_controller_001_reset_out_reset), // reset_out.reset_n
		.avalonmm_write_slave_writedata   (pd_fifo_in_writedata),                //        in.writedata
		.avalonmm_write_slave_write       (pd_fifo_in_write),                    //          .write
		.avalonmm_write_slave_waitrequest (pd_fifo_in_waitrequest),              //          .waitrequest
		.avalonmm_read_slave_readdata     (pd_fifo_out_readdata),                //       out.readdata
		.avalonmm_read_slave_read         (pd_fifo_out_read),                    //          .read
		.avalonmm_read_slave_waitrequest  (pd_fifo_out_waitrequest),             //          .waitrequest
		.rdclk_control_slave_address      (pd_fifo_out_csr_address),             //   out_csr.address
		.rdclk_control_slave_read         (pd_fifo_out_csr_read),                //          .read
		.rdclk_control_slave_writedata    (pd_fifo_out_csr_writedata),           //          .writedata
		.rdclk_control_slave_write        (pd_fifo_out_csr_write),               //          .write
		.rdclk_control_slave_readdata     (pd_fifo_out_csr_readdata),            //          .readdata
		.wrclk_control_slave_address      (pd_fifo_in_csr_address),              //    in_csr.address
		.wrclk_control_slave_read         (pd_fifo_in_csr_read),                 //          .read
		.wrclk_control_slave_writedata    (pd_fifo_in_csr_writedata),            //          .writedata
		.wrclk_control_slave_write        (pd_fifo_in_csr_write),                //          .write
		.wrclk_control_slave_readdata     (pd_fifo_in_csr_readdata)              //          .readdata
	);

	Mk8_InlineController_CPU_CurrCTRL_SYS_USB_GPIO pd_gpio (
		.clk        (pheriphal_clk_clk),               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset), //               reset.reset_n
		.address    (pd_gpio_s1_address),              //                  s1.address
		.write_n    (pd_gpio_s1_write_n),              //                    .write_n
		.writedata  (pd_gpio_s1_writedata),            //                    .writedata
		.chipselect (pd_gpio_s1_chipselect),           //                    .chipselect
		.readdata   (pd_gpio_s1_readdata),             //                    .readdata
		.in_port    (pd_gpio_in_port),                 // external_connection.export
		.out_port   (pd_gpio_out_port)                 //                    .export
	);

	Mk8_InlineController_CPU_CurrCTRL_SYS_Reset reset_pd (
		.clk        (pheriphal_clk_clk),               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset), //               reset.reset_n
		.address    (reset_pd_s1_address),             //                  s1.address
		.write_n    (reset_pd_s1_write_n),             //                    .write_n
		.writedata  (reset_pd_s1_writedata),           //                    .writedata
		.chipselect (reset_pd_s1_chipselect),          //                    .chipselect
		.readdata   (reset_pd_s1_readdata),            //                    .readdata
		.out_port   (reset_out_export)                 // external_connection.export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~pheriphal_reset_reset_n),           // reset_in0.reset
		.clk            (pheriphal_clk_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~pd_reset_reset_n),                      // reset_in0.reset
		.clk            (pd_clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
