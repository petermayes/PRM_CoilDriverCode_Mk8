// Mk8_InlineController_CPU_Pheriphals.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module Mk8_InlineController_CPU_Pheriphals (
		input  wire [7:0]  led_gpio_external_connection_in_port,  // led_gpio_external_connection.in_port
		output wire [7:0]  led_gpio_external_connection_out_port, //                             .out_port
		input  wire [2:0]  led_gpio_s1_address,                   //                  led_gpio_s1.address
		input  wire        led_gpio_s1_write_n,                   //                             .write_n
		input  wire [31:0] led_gpio_s1_writedata,                 //                             .writedata
		input  wire        led_gpio_s1_chipselect,                //                             .chipselect
		output wire [31:0] led_gpio_s1_readdata,                  //                             .readdata
		input  wire        pheriphal_clk_clk,                     //                pheriphal_clk.clk
		input  wire        pheriphal_reset_reset_n,               //              pheriphal_reset.reset_n
		output wire [7:0]  tp_gpio_external_connection_export,    //  tp_gpio_external_connection.export
		input  wire [2:0]  tp_gpio_s1_address,                    //                   tp_gpio_s1.address
		input  wire        tp_gpio_s1_write_n,                    //                             .write_n
		input  wire [31:0] tp_gpio_s1_writedata,                  //                             .writedata
		input  wire        tp_gpio_s1_chipselect,                 //                             .chipselect
		output wire [31:0] tp_gpio_s1_readdata                    //                             .readdata
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> [LED_GPIO:reset_n, TP_GPIO:reset_n]

	Mk8_InlineController_CPU_Pheriphals_LED_GPIO led_gpio (
		.clk        (pheriphal_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (led_gpio_s1_address),                   //                  s1.address
		.write_n    (led_gpio_s1_write_n),                   //                    .write_n
		.writedata  (led_gpio_s1_writedata),                 //                    .writedata
		.chipselect (led_gpio_s1_chipselect),                //                    .chipselect
		.readdata   (led_gpio_s1_readdata),                  //                    .readdata
		.in_port    (led_gpio_external_connection_in_port),  // external_connection.export
		.out_port   (led_gpio_external_connection_out_port)  //                    .export
	);

	Mk8_InlineController_CPU_Pheriphals_TP_GPIO tp_gpio (
		.clk        (pheriphal_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (tp_gpio_s1_address),                 //                  s1.address
		.write_n    (tp_gpio_s1_write_n),                 //                    .write_n
		.writedata  (tp_gpio_s1_writedata),               //                    .writedata
		.chipselect (tp_gpio_s1_chipselect),              //                    .chipselect
		.readdata   (tp_gpio_s1_readdata),                //                    .readdata
		.out_port   (tp_gpio_external_connection_export)  // external_connection.export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~pheriphal_reset_reset_n),       // reset_in0.reset
		.clk            (pheriphal_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
