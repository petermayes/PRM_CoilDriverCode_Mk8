// Mk8_InlineController_CPU.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module Mk8_InlineController_CPU (
		output wire        altpll_sys_locked_conduit_export,                 //               altpll_sys_locked_conduit.export
		input  wire        clk_clk,                                          //                                     clk.clk
		output wire        clk_10m_clk,                                      //                                 clk_10m.clk
		input  wire        clk_currctrl_fifo_clk,                            //                       clk_currctrl_fifo.clk
		input  wire        clk_currctrl_ram_clk,                             //                        clk_currctrl_ram.clk
		input  wire        clk_parameter_ram_clk_clk,                        //                   clk_parameter_ram_clk.clk
		input  wire        clk_usb_ext_clk_clk,                              //                         clk_usb_ext_clk.clk
		output wire        cpu_clk_clk,                                      //                                 cpu_clk.clk
		input  wire        currctrl_sys_bridge_acknowledge,                  //                     currctrl_sys_bridge.acknowledge
		input  wire        currctrl_sys_bridge_irq,                          //                                        .irq
		output wire [6:0]  currctrl_sys_bridge_address,                      //                                        .address
		output wire        currctrl_sys_bridge_bus_enable,                   //                                        .bus_enable
		output wire [3:0]  currctrl_sys_bridge_byte_enable,                  //                                        .byte_enable
		output wire        currctrl_sys_bridge_rw,                           //                                        .rw
		output wire [31:0] currctrl_sys_bridge_write_data,                   //                                        .write_data
		input  wire [31:0] currctrl_sys_bridge_read_data,                    //                                        .read_data
		input  wire [31:0] currctrl_sys_currctrl_gpio_ext_in_port,           //          currctrl_sys_currctrl_gpio_ext.in_port
		output wire [31:0] currctrl_sys_currctrl_gpio_ext_out_port,          //                                        .out_port
		input  wire [7:0]  currctrl_sys_register_ram_s2_address,             //            currctrl_sys_register_ram_s2.address
		input  wire        currctrl_sys_register_ram_s2_chipselect,          //                                        .chipselect
		input  wire        currctrl_sys_register_ram_s2_clken,               //                                        .clken
		input  wire        currctrl_sys_register_ram_s2_write,               //                                        .write
		output wire [31:0] currctrl_sys_register_ram_s2_readdata,            //                                        .readdata
		input  wire [31:0] currctrl_sys_register_ram_s2_writedata,           //                                        .writedata
		input  wire [3:0]  currctrl_sys_register_ram_s2_byteenable,          //                                        .byteenable
		input  wire        parameter_sys_crc_init_bridge_acknowledge,        //           parameter_sys_crc_init_bridge.acknowledge
		input  wire        parameter_sys_crc_init_bridge_irq,                //                                        .irq
		output wire [7:0]  parameter_sys_crc_init_bridge_address,            //                                        .address
		output wire        parameter_sys_crc_init_bridge_bus_enable,         //                                        .bus_enable
		output wire        parameter_sys_crc_init_bridge_byte_enable,        //                                        .byte_enable
		output wire        parameter_sys_crc_init_bridge_rw,                 //                                        .rw
		output wire [7:0]  parameter_sys_crc_init_bridge_write_data,         //                                        .write_data
		input  wire [7:0]  parameter_sys_crc_init_bridge_read_data,          //                                        .read_data
		input  wire        parameter_sys_parameter_gpio_in_port,             //            parameter_sys_parameter_gpio.in_port
		output wire        parameter_sys_parameter_gpio_out_port,            //                                        .out_port
		input  wire [10:0] parameter_sys_parameter_rx_ram_s2_address,        //       parameter_sys_parameter_rx_ram_s2.address
		input  wire        parameter_sys_parameter_rx_ram_s2_chipselect,     //                                        .chipselect
		input  wire        parameter_sys_parameter_rx_ram_s2_clken,          //                                        .clken
		input  wire        parameter_sys_parameter_rx_ram_s2_write,          //                                        .write
		output wire [31:0] parameter_sys_parameter_rx_ram_s2_readdata,       //                                        .readdata
		input  wire [31:0] parameter_sys_parameter_rx_ram_s2_writedata,      //                                        .writedata
		input  wire [3:0]  parameter_sys_parameter_rx_ram_s2_byteenable,     //                                        .byteenable
		input  wire [10:0] parameter_sys_parameter_tx_ram_s2_address,        //       parameter_sys_parameter_tx_ram_s2.address
		input  wire        parameter_sys_parameter_tx_ram_s2_chipselect,     //                                        .chipselect
		input  wire        parameter_sys_parameter_tx_ram_s2_clken,          //                                        .clken
		input  wire        parameter_sys_parameter_tx_ram_s2_write,          //                                        .write
		output wire [31:0] parameter_sys_parameter_tx_ram_s2_readdata,       //                                        .readdata
		input  wire [31:0] parameter_sys_parameter_tx_ram_s2_writedata,      //                                        .writedata
		input  wire [3:0]  parameter_sys_parameter_tx_ram_s2_byteenable,     //                                        .byteenable
		output wire [15:0] parameter_sys_parameterlengthpage_export,         //       parameter_sys_parameterlengthpage.export
		input  wire [7:0]  pheriphals_led_gpio_external_connection_in_port,  // pheriphals_led_gpio_external_connection.in_port
		output wire [7:0]  pheriphals_led_gpio_external_connection_out_port, //                                        .out_port
		output wire [7:0]  pheriphals_tp_gpio_external_connection_export,    //  pheriphals_tp_gpio_external_connection.export
		input  wire        reset_reset_n,                                    //                                   reset.reset_n
		input  wire        reset_currctrl_fifo_reset_n,                      //                     reset_currctrl_fifo.reset_n
		input  wire        reset_currctrl_ram_reset_n,                       //                      reset_currctrl_ram.reset_n
		input  wire        reset_parameter_ram_clk_reset_n,                  //                 reset_parameter_ram_clk.reset_n
		input  wire        reset_usb_ext_clk_reset_n,                        //                       reset_usb_ext_clk.reset_n
		input  wire        usb_data_sys_usb_data_gpio_in_port,               //              usb_data_sys_usb_data_gpio.in_port
		output wire        usb_data_sys_usb_data_gpio_out_port,              //                                        .out_port
		input  wire [10:0] usb_data_sys_usb_data_ram_s2_address,             //            usb_data_sys_usb_data_ram_s2.address
		input  wire        usb_data_sys_usb_data_ram_s2_chipselect,          //                                        .chipselect
		input  wire        usb_data_sys_usb_data_ram_s2_clken,               //                                        .clken
		input  wire        usb_data_sys_usb_data_ram_s2_write,               //                                        .write
		output wire [31:0] usb_data_sys_usb_data_ram_s2_readdata,            //                                        .readdata
		input  wire [31:0] usb_data_sys_usb_data_ram_s2_writedata,           //                                        .writedata
		input  wire [3:0]  usb_data_sys_usb_data_ram_s2_byteenable           //                                        .byteenable
	);

	wire          vic_0_interrupt_controller_out_valid;                                             // vic_0:interrupt_controller_out_valid -> nios2_gen2:eic_port_valid
	wire   [44:0] vic_0_interrupt_controller_out_data;                                              // vic_0:interrupt_controller_out_data -> nios2_gen2:eic_port_data
	wire          altpll_sys_c0_clk;                                                                // altpll_sys:c0 -> [CurrCTRL_SYS:cpu_clk_clk, Data_Memory:clk, Parameter_SYS:cpu_clk_clk, Program_Memory:clk, USB_Data_SYS:cpu_clk_clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, irq_synchronizer_004:sender_clk, irq_synchronizer_005:sender_clk, irq_synchronizer_006:sender_clk, mm_clock_crossing_bridge_1:s0_clk, mm_interconnect_0:altpll_sys_c0_clk, msgdma_0:clock_clk, nios2_gen2:clk, rst_controller:clk, rst_controller_002:clk, vic_0:clk_clk]
	wire          nios2_gen2_custom_instruction_master_readra;                                      // nios2_gen2:E_ci_combo_readra -> nios2_gen2_custom_instruction_master_translator:ci_slave_readra
	wire          nios2_gen2_custom_instruction_master_readrb;                                      // nios2_gen2:E_ci_combo_readrb -> nios2_gen2_custom_instruction_master_translator:ci_slave_readrb
	wire    [4:0] nios2_gen2_custom_instruction_master_multi_b;                                     // nios2_gen2:A_ci_multi_b -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_b
	wire    [4:0] nios2_gen2_custom_instruction_master_multi_c;                                     // nios2_gen2:A_ci_multi_c -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_c
	wire          nios2_gen2_custom_instruction_master_reset_req;                                   // nios2_gen2:A_ci_multi_reset_req -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire    [4:0] nios2_gen2_custom_instruction_master_multi_a;                                     // nios2_gen2:A_ci_multi_a -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_a
	wire   [31:0] nios2_gen2_custom_instruction_master_result;                                      // nios2_gen2_custom_instruction_master_translator:ci_slave_result -> nios2_gen2:E_ci_combo_result
	wire   [31:0] nios2_gen2_custom_instruction_master_datab;                                       // nios2_gen2:E_ci_combo_datab -> nios2_gen2_custom_instruction_master_translator:ci_slave_datab
	wire   [31:0] nios2_gen2_custom_instruction_master_dataa;                                       // nios2_gen2:E_ci_combo_dataa -> nios2_gen2_custom_instruction_master_translator:ci_slave_dataa
	wire          nios2_gen2_custom_instruction_master_writerc;                                     // nios2_gen2:E_ci_combo_writerc -> nios2_gen2_custom_instruction_master_translator:ci_slave_writerc
	wire   [31:0] nios2_gen2_custom_instruction_master_multi_dataa;                                 // nios2_gen2:A_ci_multi_dataa -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_dataa
	wire          nios2_gen2_custom_instruction_master_multi_writerc;                               // nios2_gen2:A_ci_multi_writerc -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_writerc
	wire    [4:0] nios2_gen2_custom_instruction_master_a;                                           // nios2_gen2:E_ci_combo_a -> nios2_gen2_custom_instruction_master_translator:ci_slave_a
	wire    [4:0] nios2_gen2_custom_instruction_master_b;                                           // nios2_gen2:E_ci_combo_b -> nios2_gen2_custom_instruction_master_translator:ci_slave_b
	wire   [31:0] nios2_gen2_custom_instruction_master_multi_result;                                // nios2_gen2_custom_instruction_master_translator:ci_slave_multi_result -> nios2_gen2:A_ci_multi_result
	wire          nios2_gen2_custom_instruction_master_clk;                                         // nios2_gen2:A_ci_multi_clock -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_clk
	wire   [31:0] nios2_gen2_custom_instruction_master_multi_datab;                                 // nios2_gen2:A_ci_multi_datab -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_datab
	wire    [4:0] nios2_gen2_custom_instruction_master_c;                                           // nios2_gen2:E_ci_combo_c -> nios2_gen2_custom_instruction_master_translator:ci_slave_c
	wire   [31:0] nios2_gen2_custom_instruction_master_ipending;                                    // nios2_gen2:E_ci_combo_ipending -> nios2_gen2_custom_instruction_master_translator:ci_slave_ipending
	wire          nios2_gen2_custom_instruction_master_start;                                       // nios2_gen2:A_ci_multi_start -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_start
	wire          nios2_gen2_custom_instruction_master_done;                                        // nios2_gen2_custom_instruction_master_translator:ci_slave_multi_done -> nios2_gen2:A_ci_multi_done
	wire    [7:0] nios2_gen2_custom_instruction_master_n;                                           // nios2_gen2:E_ci_combo_n -> nios2_gen2_custom_instruction_master_translator:ci_slave_n
	wire          nios2_gen2_custom_instruction_master_estatus;                                     // nios2_gen2:E_ci_combo_estatus -> nios2_gen2_custom_instruction_master_translator:ci_slave_estatus
	wire          nios2_gen2_custom_instruction_master_clk_en;                                      // nios2_gen2:A_ci_multi_clk_en -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_clken
	wire          nios2_gen2_custom_instruction_master_reset;                                       // nios2_gen2:A_ci_multi_reset -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_reset
	wire          nios2_gen2_custom_instruction_master_multi_readrb;                                // nios2_gen2:A_ci_multi_readrb -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_readrb
	wire          nios2_gen2_custom_instruction_master_multi_readra;                                // nios2_gen2:A_ci_multi_readra -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_readra
	wire    [7:0] nios2_gen2_custom_instruction_master_multi_n;                                     // nios2_gen2:A_ci_multi_n -> nios2_gen2_custom_instruction_master_translator:ci_slave_multi_n
	wire   [31:0] nios2_gen2_custom_instruction_master_translator_comb_ci_master_result;            // nios2_gen2_custom_instruction_master_comb_xconnect:ci_slave_result -> nios2_gen2_custom_instruction_master_translator:comb_ci_master_result
	wire          nios2_gen2_custom_instruction_master_translator_comb_ci_master_readra;            // nios2_gen2_custom_instruction_master_translator:comb_ci_master_readra -> nios2_gen2_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire    [4:0] nios2_gen2_custom_instruction_master_translator_comb_ci_master_a;                 // nios2_gen2_custom_instruction_master_translator:comb_ci_master_a -> nios2_gen2_custom_instruction_master_comb_xconnect:ci_slave_a
	wire    [4:0] nios2_gen2_custom_instruction_master_translator_comb_ci_master_b;                 // nios2_gen2_custom_instruction_master_translator:comb_ci_master_b -> nios2_gen2_custom_instruction_master_comb_xconnect:ci_slave_b
	wire          nios2_gen2_custom_instruction_master_translator_comb_ci_master_readrb;            // nios2_gen2_custom_instruction_master_translator:comb_ci_master_readrb -> nios2_gen2_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire    [4:0] nios2_gen2_custom_instruction_master_translator_comb_ci_master_c;                 // nios2_gen2_custom_instruction_master_translator:comb_ci_master_c -> nios2_gen2_custom_instruction_master_comb_xconnect:ci_slave_c
	wire          nios2_gen2_custom_instruction_master_translator_comb_ci_master_estatus;           // nios2_gen2_custom_instruction_master_translator:comb_ci_master_estatus -> nios2_gen2_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire   [31:0] nios2_gen2_custom_instruction_master_translator_comb_ci_master_ipending;          // nios2_gen2_custom_instruction_master_translator:comb_ci_master_ipending -> nios2_gen2_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire   [31:0] nios2_gen2_custom_instruction_master_translator_comb_ci_master_datab;             // nios2_gen2_custom_instruction_master_translator:comb_ci_master_datab -> nios2_gen2_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire   [31:0] nios2_gen2_custom_instruction_master_translator_comb_ci_master_dataa;             // nios2_gen2_custom_instruction_master_translator:comb_ci_master_dataa -> nios2_gen2_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire          nios2_gen2_custom_instruction_master_translator_comb_ci_master_writerc;           // nios2_gen2_custom_instruction_master_translator:comb_ci_master_writerc -> nios2_gen2_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire    [7:0] nios2_gen2_custom_instruction_master_translator_comb_ci_master_n;                 // nios2_gen2_custom_instruction_master_translator:comb_ci_master_n -> nios2_gen2_custom_instruction_master_comb_xconnect:ci_slave_n
	wire   [31:0] nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_result;             // nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios2_gen2_custom_instruction_master_comb_xconnect:ci_master0_result
	wire          nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_readra;             // nios2_gen2_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire    [4:0] nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_a;                  // nios2_gen2_custom_instruction_master_comb_xconnect:ci_master0_a -> nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire    [4:0] nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_b;                  // nios2_gen2_custom_instruction_master_comb_xconnect:ci_master0_b -> nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire          nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_readrb;             // nios2_gen2_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire    [4:0] nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_c;                  // nios2_gen2_custom_instruction_master_comb_xconnect:ci_master0_c -> nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire          nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_estatus;            // nios2_gen2_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire   [31:0] nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_ipending;           // nios2_gen2_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire   [31:0] nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_datab;              // nios2_gen2_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire   [31:0] nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_dataa;              // nios2_gen2_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire          nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_writerc;            // nios2_gen2_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire    [7:0] nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_n;                  // nios2_gen2_custom_instruction_master_comb_xconnect:ci_master0_n -> nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire   [31:0] nios2_gen2_custom_instruction_master_comb_slave_translator0_ci_master_result;     // nios_custom_instr_floating_point_2_0:s1_result -> nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire   [31:0] nios2_gen2_custom_instruction_master_comb_slave_translator0_ci_master_datab;      // nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s1_datab
	wire   [31:0] nios2_gen2_custom_instruction_master_comb_slave_translator0_ci_master_dataa;      // nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s1_dataa
	wire    [3:0] nios2_gen2_custom_instruction_master_comb_slave_translator0_ci_master_n;          // nios2_gen2_custom_instruction_master_comb_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s1_n
	wire          nios2_gen2_custom_instruction_master_translator_multi_ci_master_readra;           // nios2_gen2_custom_instruction_master_translator:multi_ci_master_readra -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire    [4:0] nios2_gen2_custom_instruction_master_translator_multi_ci_master_a;                // nios2_gen2_custom_instruction_master_translator:multi_ci_master_a -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_a
	wire    [4:0] nios2_gen2_custom_instruction_master_translator_multi_ci_master_b;                // nios2_gen2_custom_instruction_master_translator:multi_ci_master_b -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_b
	wire          nios2_gen2_custom_instruction_master_translator_multi_ci_master_clk;              // nios2_gen2_custom_instruction_master_translator:multi_ci_master_clk -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire          nios2_gen2_custom_instruction_master_translator_multi_ci_master_readrb;           // nios2_gen2_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire    [4:0] nios2_gen2_custom_instruction_master_translator_multi_ci_master_c;                // nios2_gen2_custom_instruction_master_translator:multi_ci_master_c -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_c
	wire          nios2_gen2_custom_instruction_master_translator_multi_ci_master_start;            // nios2_gen2_custom_instruction_master_translator:multi_ci_master_start -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_start
	wire          nios2_gen2_custom_instruction_master_translator_multi_ci_master_reset_req;        // nios2_gen2_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire          nios2_gen2_custom_instruction_master_translator_multi_ci_master_done;             // nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_gen2_custom_instruction_master_translator:multi_ci_master_done
	wire    [7:0] nios2_gen2_custom_instruction_master_translator_multi_ci_master_n;                // nios2_gen2_custom_instruction_master_translator:multi_ci_master_n -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_n
	wire   [31:0] nios2_gen2_custom_instruction_master_translator_multi_ci_master_result;           // nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_gen2_custom_instruction_master_translator:multi_ci_master_result
	wire          nios2_gen2_custom_instruction_master_translator_multi_ci_master_clk_en;           // nios2_gen2_custom_instruction_master_translator:multi_ci_master_clken -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire   [31:0] nios2_gen2_custom_instruction_master_translator_multi_ci_master_datab;            // nios2_gen2_custom_instruction_master_translator:multi_ci_master_datab -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire   [31:0] nios2_gen2_custom_instruction_master_translator_multi_ci_master_dataa;            // nios2_gen2_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire          nios2_gen2_custom_instruction_master_translator_multi_ci_master_reset;            // nios2_gen2_custom_instruction_master_translator:multi_ci_master_reset -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire          nios2_gen2_custom_instruction_master_translator_multi_ci_master_writerc;          // nios2_gen2_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire          nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_readra;            // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire    [4:0] nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_a;                 // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire    [4:0] nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_b;                 // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire          nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_readrb;            // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire    [4:0] nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_c;                 // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire          nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_clk;               // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire   [31:0] nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_ipending;          // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire          nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_start;             // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire          nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_reset_req;         // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire          nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_done;              // nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_done
	wire    [7:0] nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_n;                 // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire   [31:0] nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_result;            // nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_result
	wire          nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_estatus;           // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire          nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_clk_en;            // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [31:0] nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_datab;             // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire   [31:0] nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_dataa;             // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire          nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_reset;             // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire          nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_writerc;           // nios2_gen2_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire   [31:0] nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_result;    // nios_custom_instr_floating_point_2_0:s2_result -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire          nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_clk;       // nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_master_clk -> nios_custom_instr_floating_point_2_0:s2_clk
	wire          nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;    // nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_master_clken -> nios_custom_instr_floating_point_2_0:s2_clk_en
	wire   [31:0] nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_datab;     // nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s2_datab
	wire   [31:0] nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_dataa;     // nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s2_dataa
	wire          nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_start;     // nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_master_start -> nios_custom_instr_floating_point_2_0:s2_start
	wire          nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_reset;     // nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_master_reset -> nios_custom_instr_floating_point_2_0:s2_reset
	wire          nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_reset_req; // nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> nios_custom_instr_floating_point_2_0:s2_reset_req
	wire          nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_done;      // nios_custom_instr_floating_point_2_0:s2_done -> nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire    [2:0] nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_n;         // nios2_gen2_custom_instruction_master_multi_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s2_n
	wire   [31:0] nios2_gen2_data_master_readdata;                                                  // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire          nios2_gen2_data_master_waitrequest;                                               // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire          nios2_gen2_data_master_debugaccess;                                               // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire   [25:0] nios2_gen2_data_master_address;                                                   // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire    [3:0] nios2_gen2_data_master_byteenable;                                                // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire          nios2_gen2_data_master_read;                                                      // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire          nios2_gen2_data_master_write;                                                     // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire   [31:0] nios2_gen2_data_master_writedata;                                                 // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire   [31:0] msgdma_0_mm_read_readdata;                                                        // mm_interconnect_0:msgdma_0_mm_read_readdata -> msgdma_0:mm_read_readdata
	wire          msgdma_0_mm_read_waitrequest;                                                     // mm_interconnect_0:msgdma_0_mm_read_waitrequest -> msgdma_0:mm_read_waitrequest
	wire   [24:0] msgdma_0_mm_read_address;                                                         // msgdma_0:mm_read_address -> mm_interconnect_0:msgdma_0_mm_read_address
	wire          msgdma_0_mm_read_read;                                                            // msgdma_0:mm_read_read -> mm_interconnect_0:msgdma_0_mm_read_read
	wire    [3:0] msgdma_0_mm_read_byteenable;                                                      // msgdma_0:mm_read_byteenable -> mm_interconnect_0:msgdma_0_mm_read_byteenable
	wire          msgdma_0_mm_read_readdatavalid;                                                   // mm_interconnect_0:msgdma_0_mm_read_readdatavalid -> msgdma_0:mm_read_readdatavalid
	wire          msgdma_0_mm_write_waitrequest;                                                    // mm_interconnect_0:msgdma_0_mm_write_waitrequest -> msgdma_0:mm_write_waitrequest
	wire   [24:0] msgdma_0_mm_write_address;                                                        // msgdma_0:mm_write_address -> mm_interconnect_0:msgdma_0_mm_write_address
	wire    [3:0] msgdma_0_mm_write_byteenable;                                                     // msgdma_0:mm_write_byteenable -> mm_interconnect_0:msgdma_0_mm_write_byteenable
	wire          msgdma_0_mm_write_write;                                                          // msgdma_0:mm_write_write -> mm_interconnect_0:msgdma_0_mm_write_write
	wire   [31:0] msgdma_0_mm_write_writedata;                                                      // msgdma_0:mm_write_writedata -> mm_interconnect_0:msgdma_0_mm_write_writedata
	wire   [31:0] nios2_gen2_instruction_master_readdata;                                           // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire          nios2_gen2_instruction_master_waitrequest;                                        // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire   [16:0] nios2_gen2_instruction_master_address;                                            // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire          nios2_gen2_instruction_master_read;                                               // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire          nios2_gen2_instruction_master_readdatavalid;                                      // mm_interconnect_0:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire   [31:0] mm_interconnect_0_msgdma_0_csr_readdata;                                          // msgdma_0:csr_readdata -> mm_interconnect_0:msgdma_0_csr_readdata
	wire    [2:0] mm_interconnect_0_msgdma_0_csr_address;                                           // mm_interconnect_0:msgdma_0_csr_address -> msgdma_0:csr_address
	wire          mm_interconnect_0_msgdma_0_csr_read;                                              // mm_interconnect_0:msgdma_0_csr_read -> msgdma_0:csr_read
	wire    [3:0] mm_interconnect_0_msgdma_0_csr_byteenable;                                        // mm_interconnect_0:msgdma_0_csr_byteenable -> msgdma_0:csr_byteenable
	wire          mm_interconnect_0_msgdma_0_csr_write;                                             // mm_interconnect_0:msgdma_0_csr_write -> msgdma_0:csr_write
	wire   [31:0] mm_interconnect_0_msgdma_0_csr_writedata;                                         // mm_interconnect_0:msgdma_0_csr_writedata -> msgdma_0:csr_writedata
	wire   [31:0] mm_interconnect_0_vic_0_csr_access_readdata;                                      // vic_0:csr_access_readdata -> mm_interconnect_0:vic_0_csr_access_readdata
	wire    [7:0] mm_interconnect_0_vic_0_csr_access_address;                                       // mm_interconnect_0:vic_0_csr_access_address -> vic_0:csr_access_address
	wire          mm_interconnect_0_vic_0_csr_access_read;                                          // mm_interconnect_0:vic_0_csr_access_read -> vic_0:csr_access_read
	wire          mm_interconnect_0_vic_0_csr_access_write;                                         // mm_interconnect_0:vic_0_csr_access_write -> vic_0:csr_access_write
	wire   [31:0] mm_interconnect_0_vic_0_csr_access_writedata;                                     // mm_interconnect_0:vic_0_csr_access_writedata -> vic_0:csr_access_writedata
	wire   [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;                            // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire          mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;                         // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;                         // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;                             // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire          mm_interconnect_0_nios2_gen2_debug_mem_slave_read;                                // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;                          // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire          mm_interconnect_0_nios2_gen2_debug_mem_slave_write;                               // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;                           // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire          mm_interconnect_0_msgdma_0_descriptor_slave_waitrequest;                          // msgdma_0:descriptor_slave_waitrequest -> mm_interconnect_0:msgdma_0_descriptor_slave_waitrequest
	wire   [31:0] mm_interconnect_0_msgdma_0_descriptor_slave_byteenable;                           // mm_interconnect_0:msgdma_0_descriptor_slave_byteenable -> msgdma_0:descriptor_slave_byteenable
	wire          mm_interconnect_0_msgdma_0_descriptor_slave_write;                                // mm_interconnect_0:msgdma_0_descriptor_slave_write -> msgdma_0:descriptor_slave_write
	wire  [255:0] mm_interconnect_0_msgdma_0_descriptor_slave_writedata;                            // mm_interconnect_0:msgdma_0_descriptor_slave_writedata -> msgdma_0:descriptor_slave_writedata
	wire          mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_chipselect;                   // mm_interconnect_0:Parameter_SYS_parameter_rx_ram_s1_chipselect -> Parameter_SYS:parameter_rx_ram_s1_chipselect
	wire   [31:0] mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_readdata;                     // Parameter_SYS:parameter_rx_ram_s1_readdata -> mm_interconnect_0:Parameter_SYS_parameter_rx_ram_s1_readdata
	wire   [10:0] mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_address;                      // mm_interconnect_0:Parameter_SYS_parameter_rx_ram_s1_address -> Parameter_SYS:parameter_rx_ram_s1_address
	wire    [3:0] mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_byteenable;                   // mm_interconnect_0:Parameter_SYS_parameter_rx_ram_s1_byteenable -> Parameter_SYS:parameter_rx_ram_s1_byteenable
	wire          mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_write;                        // mm_interconnect_0:Parameter_SYS_parameter_rx_ram_s1_write -> Parameter_SYS:parameter_rx_ram_s1_write
	wire   [31:0] mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_writedata;                    // mm_interconnect_0:Parameter_SYS_parameter_rx_ram_s1_writedata -> Parameter_SYS:parameter_rx_ram_s1_writedata
	wire          mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_clken;                        // mm_interconnect_0:Parameter_SYS_parameter_rx_ram_s1_clken -> Parameter_SYS:parameter_rx_ram_s1_clken
	wire          mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_chipselect;                   // mm_interconnect_0:Parameter_SYS_parameter_tx_ram_s1_chipselect -> Parameter_SYS:parameter_tx_ram_s1_chipselect
	wire   [31:0] mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_readdata;                     // Parameter_SYS:parameter_tx_ram_s1_readdata -> mm_interconnect_0:Parameter_SYS_parameter_tx_ram_s1_readdata
	wire   [10:0] mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_address;                      // mm_interconnect_0:Parameter_SYS_parameter_tx_ram_s1_address -> Parameter_SYS:parameter_tx_ram_s1_address
	wire    [3:0] mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_byteenable;                   // mm_interconnect_0:Parameter_SYS_parameter_tx_ram_s1_byteenable -> Parameter_SYS:parameter_tx_ram_s1_byteenable
	wire          mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_write;                        // mm_interconnect_0:Parameter_SYS_parameter_tx_ram_s1_write -> Parameter_SYS:parameter_tx_ram_s1_write
	wire   [31:0] mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_writedata;                    // mm_interconnect_0:Parameter_SYS_parameter_tx_ram_s1_writedata -> Parameter_SYS:parameter_tx_ram_s1_writedata
	wire          mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_clken;                        // mm_interconnect_0:Parameter_SYS_parameter_tx_ram_s1_clken -> Parameter_SYS:parameter_tx_ram_s1_clken
	wire   [31:0] mm_interconnect_0_altpll_sys_pll_slave_readdata;                                  // altpll_sys:readdata -> mm_interconnect_0:altpll_sys_pll_slave_readdata
	wire    [1:0] mm_interconnect_0_altpll_sys_pll_slave_address;                                   // mm_interconnect_0:altpll_sys_pll_slave_address -> altpll_sys:address
	wire          mm_interconnect_0_altpll_sys_pll_slave_read;                                      // mm_interconnect_0:altpll_sys_pll_slave_read -> altpll_sys:read
	wire          mm_interconnect_0_altpll_sys_pll_slave_write;                                     // mm_interconnect_0:altpll_sys_pll_slave_write -> altpll_sys:write
	wire   [31:0] mm_interconnect_0_altpll_sys_pll_slave_writedata;                                 // mm_interconnect_0:altpll_sys_pll_slave_writedata -> altpll_sys:writedata
	wire   [31:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdata;                         // mm_clock_crossing_bridge_1:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_1_s0_readdata
	wire          mm_interconnect_0_mm_clock_crossing_bridge_1_s0_waitrequest;                      // mm_clock_crossing_bridge_1:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_1_s0_waitrequest
	wire          mm_interconnect_0_mm_clock_crossing_bridge_1_s0_debugaccess;                      // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_debugaccess -> mm_clock_crossing_bridge_1:s0_debugaccess
	wire   [10:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_address;                          // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_address -> mm_clock_crossing_bridge_1:s0_address
	wire          mm_interconnect_0_mm_clock_crossing_bridge_1_s0_read;                             // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_read -> mm_clock_crossing_bridge_1:s0_read
	wire    [3:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_byteenable;                       // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_byteenable -> mm_clock_crossing_bridge_1:s0_byteenable
	wire          mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdatavalid;                    // mm_clock_crossing_bridge_1:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_1_s0_readdatavalid
	wire          mm_interconnect_0_mm_clock_crossing_bridge_1_s0_write;                            // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_write -> mm_clock_crossing_bridge_1:s0_write
	wire   [31:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_writedata;                        // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_writedata -> mm_clock_crossing_bridge_1:s0_writedata
	wire    [0:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_burstcount;                       // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_burstcount -> mm_clock_crossing_bridge_1:s0_burstcount
	wire          mm_interconnect_0_program_memory_s1_chipselect;                                   // mm_interconnect_0:Program_Memory_s1_chipselect -> Program_Memory:chipselect
	wire   [31:0] mm_interconnect_0_program_memory_s1_readdata;                                     // Program_Memory:readdata -> mm_interconnect_0:Program_Memory_s1_readdata
	wire   [12:0] mm_interconnect_0_program_memory_s1_address;                                      // mm_interconnect_0:Program_Memory_s1_address -> Program_Memory:address
	wire    [3:0] mm_interconnect_0_program_memory_s1_byteenable;                                   // mm_interconnect_0:Program_Memory_s1_byteenable -> Program_Memory:byteenable
	wire          mm_interconnect_0_program_memory_s1_write;                                        // mm_interconnect_0:Program_Memory_s1_write -> Program_Memory:write
	wire   [31:0] mm_interconnect_0_program_memory_s1_writedata;                                    // mm_interconnect_0:Program_Memory_s1_writedata -> Program_Memory:writedata
	wire          mm_interconnect_0_program_memory_s1_clken;                                        // mm_interconnect_0:Program_Memory_s1_clken -> Program_Memory:clken
	wire          mm_interconnect_0_data_memory_s1_chipselect;                                      // mm_interconnect_0:Data_Memory_s1_chipselect -> Data_Memory:chipselect
	wire   [31:0] mm_interconnect_0_data_memory_s1_readdata;                                        // Data_Memory:readdata -> mm_interconnect_0:Data_Memory_s1_readdata
	wire   [11:0] mm_interconnect_0_data_memory_s1_address;                                         // mm_interconnect_0:Data_Memory_s1_address -> Data_Memory:address
	wire    [3:0] mm_interconnect_0_data_memory_s1_byteenable;                                      // mm_interconnect_0:Data_Memory_s1_byteenable -> Data_Memory:byteenable
	wire          mm_interconnect_0_data_memory_s1_write;                                           // mm_interconnect_0:Data_Memory_s1_write -> Data_Memory:write
	wire   [31:0] mm_interconnect_0_data_memory_s1_writedata;                                       // mm_interconnect_0:Data_Memory_s1_writedata -> Data_Memory:writedata
	wire          mm_interconnect_0_data_memory_s1_clken;                                           // mm_interconnect_0:Data_Memory_s1_clken -> Data_Memory:clken
	wire          mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_chipselect;                          // mm_interconnect_0:USB_Data_SYS_usb_rx_ram_s1_chipselect -> USB_Data_SYS:usb_rx_ram_s1_chipselect
	wire   [31:0] mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_readdata;                            // USB_Data_SYS:usb_rx_ram_s1_readdata -> mm_interconnect_0:USB_Data_SYS_usb_rx_ram_s1_readdata
	wire   [10:0] mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_address;                             // mm_interconnect_0:USB_Data_SYS_usb_rx_ram_s1_address -> USB_Data_SYS:usb_rx_ram_s1_address
	wire    [3:0] mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_byteenable;                          // mm_interconnect_0:USB_Data_SYS_usb_rx_ram_s1_byteenable -> USB_Data_SYS:usb_rx_ram_s1_byteenable
	wire          mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_write;                               // mm_interconnect_0:USB_Data_SYS_usb_rx_ram_s1_write -> USB_Data_SYS:usb_rx_ram_s1_write
	wire   [31:0] mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_writedata;                           // mm_interconnect_0:USB_Data_SYS_usb_rx_ram_s1_writedata -> USB_Data_SYS:usb_rx_ram_s1_writedata
	wire          mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_clken;                               // mm_interconnect_0:USB_Data_SYS_usb_rx_ram_s1_clken -> USB_Data_SYS:usb_rx_ram_s1_clken
	wire          mm_clock_crossing_bridge_1_m0_waitrequest;                                        // mm_interconnect_1:mm_clock_crossing_bridge_1_m0_waitrequest -> mm_clock_crossing_bridge_1:m0_waitrequest
	wire   [31:0] mm_clock_crossing_bridge_1_m0_readdata;                                           // mm_interconnect_1:mm_clock_crossing_bridge_1_m0_readdata -> mm_clock_crossing_bridge_1:m0_readdata
	wire          mm_clock_crossing_bridge_1_m0_debugaccess;                                        // mm_clock_crossing_bridge_1:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_debugaccess
	wire   [10:0] mm_clock_crossing_bridge_1_m0_address;                                            // mm_clock_crossing_bridge_1:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_address
	wire          mm_clock_crossing_bridge_1_m0_read;                                               // mm_clock_crossing_bridge_1:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_read
	wire    [3:0] mm_clock_crossing_bridge_1_m0_byteenable;                                         // mm_clock_crossing_bridge_1:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_byteenable
	wire          mm_clock_crossing_bridge_1_m0_readdatavalid;                                      // mm_interconnect_1:mm_clock_crossing_bridge_1_m0_readdatavalid -> mm_clock_crossing_bridge_1:m0_readdatavalid
	wire   [31:0] mm_clock_crossing_bridge_1_m0_writedata;                                          // mm_clock_crossing_bridge_1:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_writedata
	wire          mm_clock_crossing_bridge_1_m0_write;                                              // mm_clock_crossing_bridge_1:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_write
	wire    [0:0] mm_clock_crossing_bridge_1_m0_burstcount;                                         // mm_clock_crossing_bridge_1:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_burstcount
	wire          mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_chipselect;          // mm_interconnect_1:Parameter_SYS_crc_init_bridge_avalon_slave_chipselect -> Parameter_SYS:crc_init_bridge_avalon_slave_chipselect
	wire    [7:0] mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_readdata;            // Parameter_SYS:crc_init_bridge_avalon_slave_readdata -> mm_interconnect_1:Parameter_SYS_crc_init_bridge_avalon_slave_readdata
	wire          mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_waitrequest;         // Parameter_SYS:crc_init_bridge_avalon_slave_waitrequest -> mm_interconnect_1:Parameter_SYS_crc_init_bridge_avalon_slave_waitrequest
	wire    [7:0] mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_address;             // mm_interconnect_1:Parameter_SYS_crc_init_bridge_avalon_slave_address -> Parameter_SYS:crc_init_bridge_avalon_slave_address
	wire          mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_read;                // mm_interconnect_1:Parameter_SYS_crc_init_bridge_avalon_slave_read -> Parameter_SYS:crc_init_bridge_avalon_slave_read
	wire    [0:0] mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_byteenable;          // mm_interconnect_1:Parameter_SYS_crc_init_bridge_avalon_slave_byteenable -> Parameter_SYS:crc_init_bridge_avalon_slave_byteenable
	wire          mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_write;               // mm_interconnect_1:Parameter_SYS_crc_init_bridge_avalon_slave_write -> Parameter_SYS:crc_init_bridge_avalon_slave_write
	wire    [7:0] mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_writedata;           // mm_interconnect_1:Parameter_SYS_crc_init_bridge_avalon_slave_writedata -> Parameter_SYS:crc_init_bridge_avalon_slave_writedata
	wire          mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_chipselect;                       // mm_interconnect_1:CurrCTRL_SYS_currctrl_gpio_s1_chipselect -> CurrCTRL_SYS:currctrl_gpio_s1_chipselect
	wire   [31:0] mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_readdata;                         // CurrCTRL_SYS:currctrl_gpio_s1_readdata -> mm_interconnect_1:CurrCTRL_SYS_currctrl_gpio_s1_readdata
	wire    [2:0] mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_address;                          // mm_interconnect_1:CurrCTRL_SYS_currctrl_gpio_s1_address -> CurrCTRL_SYS:currctrl_gpio_s1_address
	wire          mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_write;                            // mm_interconnect_1:CurrCTRL_SYS_currctrl_gpio_s1_write -> CurrCTRL_SYS:currctrl_gpio_s1_write_n
	wire   [31:0] mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_writedata;                        // mm_interconnect_1:CurrCTRL_SYS_currctrl_gpio_s1_writedata -> CurrCTRL_SYS:currctrl_gpio_s1_writedata
	wire          mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_chipselect;               // mm_interconnect_1:CurrCTRL_SYS_currctrl_register_ram_s1_chipselect -> CurrCTRL_SYS:currctrl_register_ram_s1_chipselect
	wire   [31:0] mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_readdata;                 // CurrCTRL_SYS:currctrl_register_ram_s1_readdata -> mm_interconnect_1:CurrCTRL_SYS_currctrl_register_ram_s1_readdata
	wire    [7:0] mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_address;                  // mm_interconnect_1:CurrCTRL_SYS_currctrl_register_ram_s1_address -> CurrCTRL_SYS:currctrl_register_ram_s1_address
	wire    [3:0] mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_byteenable;               // mm_interconnect_1:CurrCTRL_SYS_currctrl_register_ram_s1_byteenable -> CurrCTRL_SYS:currctrl_register_ram_s1_byteenable
	wire          mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_write;                    // mm_interconnect_1:CurrCTRL_SYS_currctrl_register_ram_s1_write -> CurrCTRL_SYS:currctrl_register_ram_s1_write
	wire   [31:0] mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_writedata;                // mm_interconnect_1:CurrCTRL_SYS_currctrl_register_ram_s1_writedata -> CurrCTRL_SYS:currctrl_register_ram_s1_writedata
	wire          mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_clken;                    // mm_interconnect_1:CurrCTRL_SYS_currctrl_register_ram_s1_clken -> CurrCTRL_SYS:currctrl_register_ram_s1_clken
	wire          mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_chipselect;        // mm_interconnect_1:CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_chipselect -> CurrCTRL_SYS:currctrlsys_bridge_avalon_slave_chipselect
	wire   [31:0] mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_readdata;          // CurrCTRL_SYS:currctrlsys_bridge_avalon_slave_readdata -> mm_interconnect_1:CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_readdata
	wire          mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_waitrequest;       // CurrCTRL_SYS:currctrlsys_bridge_avalon_slave_waitrequest -> mm_interconnect_1:CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_waitrequest
	wire    [4:0] mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_address;           // mm_interconnect_1:CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_address -> CurrCTRL_SYS:currctrlsys_bridge_avalon_slave_address
	wire          mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_read;              // mm_interconnect_1:CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_read -> CurrCTRL_SYS:currctrlsys_bridge_avalon_slave_read
	wire    [3:0] mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_byteenable;        // mm_interconnect_1:CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_byteenable -> CurrCTRL_SYS:currctrlsys_bridge_avalon_slave_byteenable
	wire          mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_write;             // mm_interconnect_1:CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_write -> CurrCTRL_SYS:currctrlsys_bridge_avalon_slave_write
	wire   [31:0] mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_writedata;         // mm_interconnect_1:CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_writedata -> CurrCTRL_SYS:currctrlsys_bridge_avalon_slave_writedata
	wire          mm_interconnect_1_pheriphals_led_gpio_s1_chipselect;                              // mm_interconnect_1:Pheriphals_led_gpio_s1_chipselect -> Pheriphals:led_gpio_s1_chipselect
	wire   [31:0] mm_interconnect_1_pheriphals_led_gpio_s1_readdata;                                // Pheriphals:led_gpio_s1_readdata -> mm_interconnect_1:Pheriphals_led_gpio_s1_readdata
	wire    [2:0] mm_interconnect_1_pheriphals_led_gpio_s1_address;                                 // mm_interconnect_1:Pheriphals_led_gpio_s1_address -> Pheriphals:led_gpio_s1_address
	wire          mm_interconnect_1_pheriphals_led_gpio_s1_write;                                   // mm_interconnect_1:Pheriphals_led_gpio_s1_write -> Pheriphals:led_gpio_s1_write_n
	wire   [31:0] mm_interconnect_1_pheriphals_led_gpio_s1_writedata;                               // mm_interconnect_1:Pheriphals_led_gpio_s1_writedata -> Pheriphals:led_gpio_s1_writedata
	wire          mm_interconnect_1_parameter_sys_parameter_gpio_s1_chipselect;                     // mm_interconnect_1:Parameter_SYS_parameter_gpio_s1_chipselect -> Parameter_SYS:parameter_gpio_s1_chipselect
	wire   [31:0] mm_interconnect_1_parameter_sys_parameter_gpio_s1_readdata;                       // Parameter_SYS:parameter_gpio_s1_readdata -> mm_interconnect_1:Parameter_SYS_parameter_gpio_s1_readdata
	wire    [2:0] mm_interconnect_1_parameter_sys_parameter_gpio_s1_address;                        // mm_interconnect_1:Parameter_SYS_parameter_gpio_s1_address -> Parameter_SYS:parameter_gpio_s1_address
	wire          mm_interconnect_1_parameter_sys_parameter_gpio_s1_write;                          // mm_interconnect_1:Parameter_SYS_parameter_gpio_s1_write -> Parameter_SYS:parameter_gpio_s1_write_n
	wire   [31:0] mm_interconnect_1_parameter_sys_parameter_gpio_s1_writedata;                      // mm_interconnect_1:Parameter_SYS_parameter_gpio_s1_writedata -> Parameter_SYS:parameter_gpio_s1_writedata
	wire          mm_interconnect_1_parameter_sys_parameterlengthpage_s1_chipselect;                // mm_interconnect_1:Parameter_SYS_parameterlengthpage_s1_chipselect -> Parameter_SYS:parameterlengthpage_s1_chipselect
	wire   [31:0] mm_interconnect_1_parameter_sys_parameterlengthpage_s1_readdata;                  // Parameter_SYS:parameterlengthpage_s1_readdata -> mm_interconnect_1:Parameter_SYS_parameterlengthpage_s1_readdata
	wire    [1:0] mm_interconnect_1_parameter_sys_parameterlengthpage_s1_address;                   // mm_interconnect_1:Parameter_SYS_parameterlengthpage_s1_address -> Parameter_SYS:parameterlengthpage_s1_address
	wire          mm_interconnect_1_parameter_sys_parameterlengthpage_s1_write;                     // mm_interconnect_1:Parameter_SYS_parameterlengthpage_s1_write -> Parameter_SYS:parameterlengthpage_s1_write_n
	wire   [31:0] mm_interconnect_1_parameter_sys_parameterlengthpage_s1_writedata;                 // mm_interconnect_1:Parameter_SYS_parameterlengthpage_s1_writedata -> Parameter_SYS:parameterlengthpage_s1_writedata
	wire          mm_interconnect_1_timersys_timer_0_s1_chipselect;                                 // mm_interconnect_1:TimerSYS_timer_0_s1_chipselect -> TimerSYS:timer_0_s1_chipselect
	wire   [15:0] mm_interconnect_1_timersys_timer_0_s1_readdata;                                   // TimerSYS:timer_0_s1_readdata -> mm_interconnect_1:TimerSYS_timer_0_s1_readdata
	wire    [2:0] mm_interconnect_1_timersys_timer_0_s1_address;                                    // mm_interconnect_1:TimerSYS_timer_0_s1_address -> TimerSYS:timer_0_s1_address
	wire          mm_interconnect_1_timersys_timer_0_s1_write;                                      // mm_interconnect_1:TimerSYS_timer_0_s1_write -> TimerSYS:timer_0_s1_write_n
	wire   [15:0] mm_interconnect_1_timersys_timer_0_s1_writedata;                                  // mm_interconnect_1:TimerSYS_timer_0_s1_writedata -> TimerSYS:timer_0_s1_writedata
	wire          mm_interconnect_1_timersys_timer_1_s1_chipselect;                                 // mm_interconnect_1:TimerSYS_timer_1_s1_chipselect -> TimerSYS:timer_1_s1_chipselect
	wire   [15:0] mm_interconnect_1_timersys_timer_1_s1_readdata;                                   // TimerSYS:timer_1_s1_readdata -> mm_interconnect_1:TimerSYS_timer_1_s1_readdata
	wire    [2:0] mm_interconnect_1_timersys_timer_1_s1_address;                                    // mm_interconnect_1:TimerSYS_timer_1_s1_address -> TimerSYS:timer_1_s1_address
	wire          mm_interconnect_1_timersys_timer_1_s1_write;                                      // mm_interconnect_1:TimerSYS_timer_1_s1_write -> TimerSYS:timer_1_s1_write_n
	wire   [15:0] mm_interconnect_1_timersys_timer_1_s1_writedata;                                  // mm_interconnect_1:TimerSYS_timer_1_s1_writedata -> TimerSYS:timer_1_s1_writedata
	wire          mm_interconnect_1_timersys_timer_2_s1_chipselect;                                 // mm_interconnect_1:TimerSYS_timer_2_s1_chipselect -> TimerSYS:timer_2_s1_chipselect
	wire   [15:0] mm_interconnect_1_timersys_timer_2_s1_readdata;                                   // TimerSYS:timer_2_s1_readdata -> mm_interconnect_1:TimerSYS_timer_2_s1_readdata
	wire    [2:0] mm_interconnect_1_timersys_timer_2_s1_address;                                    // mm_interconnect_1:TimerSYS_timer_2_s1_address -> TimerSYS:timer_2_s1_address
	wire          mm_interconnect_1_timersys_timer_2_s1_write;                                      // mm_interconnect_1:TimerSYS_timer_2_s1_write -> TimerSYS:timer_2_s1_write_n
	wire   [15:0] mm_interconnect_1_timersys_timer_2_s1_writedata;                                  // mm_interconnect_1:TimerSYS_timer_2_s1_writedata -> TimerSYS:timer_2_s1_writedata
	wire          mm_interconnect_1_pheriphals_tp_gpio_s1_chipselect;                               // mm_interconnect_1:Pheriphals_tp_gpio_s1_chipselect -> Pheriphals:tp_gpio_s1_chipselect
	wire   [31:0] mm_interconnect_1_pheriphals_tp_gpio_s1_readdata;                                 // Pheriphals:tp_gpio_s1_readdata -> mm_interconnect_1:Pheriphals_tp_gpio_s1_readdata
	wire    [2:0] mm_interconnect_1_pheriphals_tp_gpio_s1_address;                                  // mm_interconnect_1:Pheriphals_tp_gpio_s1_address -> Pheriphals:tp_gpio_s1_address
	wire          mm_interconnect_1_pheriphals_tp_gpio_s1_write;                                    // mm_interconnect_1:Pheriphals_tp_gpio_s1_write -> Pheriphals:tp_gpio_s1_write_n
	wire   [31:0] mm_interconnect_1_pheriphals_tp_gpio_s1_writedata;                                // mm_interconnect_1:Pheriphals_tp_gpio_s1_writedata -> Pheriphals:tp_gpio_s1_writedata
	wire          mm_interconnect_1_usb_data_sys_usb_gpio_s1_chipselect;                            // mm_interconnect_1:USB_Data_SYS_usb_gpio_s1_chipselect -> USB_Data_SYS:usb_gpio_s1_chipselect
	wire   [31:0] mm_interconnect_1_usb_data_sys_usb_gpio_s1_readdata;                              // USB_Data_SYS:usb_gpio_s1_readdata -> mm_interconnect_1:USB_Data_SYS_usb_gpio_s1_readdata
	wire    [2:0] mm_interconnect_1_usb_data_sys_usb_gpio_s1_address;                               // mm_interconnect_1:USB_Data_SYS_usb_gpio_s1_address -> USB_Data_SYS:usb_gpio_s1_address
	wire          mm_interconnect_1_usb_data_sys_usb_gpio_s1_write;                                 // mm_interconnect_1:USB_Data_SYS_usb_gpio_s1_write -> USB_Data_SYS:usb_gpio_s1_write_n
	wire   [31:0] mm_interconnect_1_usb_data_sys_usb_gpio_s1_writedata;                             // mm_interconnect_1:USB_Data_SYS_usb_gpio_s1_writedata -> USB_Data_SYS:usb_gpio_s1_writedata
	wire          irq_mapper_receiver1_irq;                                                         // msgdma_0:csr_irq_irq -> irq_mapper:receiver1_irq
	wire    [9:0] vic_0_irq_input_irq;                                                              // irq_mapper:sender_irq -> vic_0:irq_input_irq
	wire          irq_mapper_receiver0_irq;                                                         // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                    // Parameter_SYS:crc_init_bridge_interrupt_irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver2_irq;                                                         // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                                // CurrCTRL_SYS:currctrlsys_bridge_interrupt_irq -> irq_synchronizer_001:receiver_irq
	wire          irq_mapper_receiver3_irq;                                                         // irq_synchronizer_002:sender_irq -> irq_mapper:receiver3_irq
	wire    [0:0] irq_synchronizer_002_receiver_irq;                                                // Parameter_SYS:parameter_loop_gpio_irq_irq -> irq_synchronizer_002:receiver_irq
	wire          irq_mapper_receiver4_irq;                                                         // irq_synchronizer_003:sender_irq -> irq_mapper:receiver4_irq
	wire    [0:0] irq_synchronizer_003_receiver_irq;                                                // TimerSYS:timer_0_irq_irq -> irq_synchronizer_003:receiver_irq
	wire          irq_mapper_receiver5_irq;                                                         // irq_synchronizer_004:sender_irq -> irq_mapper:receiver5_irq
	wire    [0:0] irq_synchronizer_004_receiver_irq;                                                // TimerSYS:timer_1_irq_irq -> irq_synchronizer_004:receiver_irq
	wire          irq_mapper_receiver6_irq;                                                         // irq_synchronizer_005:sender_irq -> irq_mapper:receiver6_irq
	wire    [0:0] irq_synchronizer_005_receiver_irq;                                                // TimerSYS:timer_2_irq_irq -> irq_synchronizer_005:receiver_irq
	wire          irq_mapper_receiver7_irq;                                                         // irq_synchronizer_006:sender_irq -> irq_mapper:receiver7_irq
	wire    [0:0] irq_synchronizer_006_receiver_irq;                                                // USB_Data_SYS:usb_data_gpio_irq_irq -> irq_synchronizer_006:receiver_irq
	wire          rst_controller_reset_out_reset;                                                   // rst_controller:reset_out -> [Data_Memory:reset, Program_Memory:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, irq_synchronizer_006:sender_reset, mm_clock_crossing_bridge_1:s0_reset, mm_interconnect_0:Parameter_SYS_cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_0:msgdma_0_reset_n_reset_bridge_in_reset_reset, msgdma_0:reset_n_reset_n, rst_translator:in_reset, vic_0:reset_reset]
	wire          rst_controller_reset_out_reset_req;                                               // rst_controller:reset_req -> [Data_Memory:reset_req, Program_Memory:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                                               // rst_controller_001:reset_out -> [altpll_sys:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, irq_synchronizer_005:receiver_reset, irq_synchronizer_006:receiver_reset, mm_clock_crossing_bridge_1:m0_reset, mm_interconnect_0:altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset, mm_interconnect_1:Parameter_SYS_pheriphal_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_clock_crossing_bridge_1_m0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                                               // rst_controller_002:reset_out -> [mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n]
	wire          rst_controller_002_reset_out_reset_req;                                           // rst_controller_002:reset_req -> nios2_gen2:reset_req
	wire          nios2_gen2_debug_reset_request_reset;                                             // nios2_gen2:debug_reset_request -> rst_controller_002:reset_in1

	Mk8_InlineController_CPU_CurrCTRL_SYS currctrl_sys (
		.clk_currctrl_sys_fifo_clk                   (clk_currctrl_fifo_clk),                                                      //           clk_currctrl_sys_fifo.clk
		.clk_currctrl_sys_ram_clk                    (clk_currctrl_ram_clk),                                                       //            clk_currctrl_sys_ram.clk
		.clk_pheripal_clk                            (clk_clk),                                                                    //                    clk_pheripal.clk
		.cpu_clk_clk                                 (altpll_sys_c0_clk),                                                          //                         cpu_clk.clk
		.cpu_reset_reset_n                           (reset_reset_n),                                                              //                       cpu_reset.reset_n
		.currctrl_gpio_ext_in_port                   (currctrl_sys_currctrl_gpio_ext_in_port),                                     //               currctrl_gpio_ext.in_port
		.currctrl_gpio_ext_out_port                  (currctrl_sys_currctrl_gpio_ext_out_port),                                    //                                .out_port
		.currctrl_gpio_s1_address                    (mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_address),                    //                currctrl_gpio_s1.address
		.currctrl_gpio_s1_write_n                    (~mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_write),                     //                                .write_n
		.currctrl_gpio_s1_writedata                  (mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_writedata),                  //                                .writedata
		.currctrl_gpio_s1_chipselect                 (mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_chipselect),                 //                                .chipselect
		.currctrl_gpio_s1_readdata                   (mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_readdata),                   //                                .readdata
		.currctrl_register_ram_s1_address            (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_address),            //        currctrl_register_ram_s1.address
		.currctrl_register_ram_s1_clken              (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_clken),              //                                .clken
		.currctrl_register_ram_s1_chipselect         (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_chipselect),         //                                .chipselect
		.currctrl_register_ram_s1_write              (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_write),              //                                .write
		.currctrl_register_ram_s1_readdata           (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_readdata),           //                                .readdata
		.currctrl_register_ram_s1_writedata          (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_writedata),          //                                .writedata
		.currctrl_register_ram_s1_byteenable         (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_byteenable),         //                                .byteenable
		.currctrl_register_ram_s2_address            (currctrl_sys_register_ram_s2_address),                                       //        currctrl_register_ram_s2.address
		.currctrl_register_ram_s2_chipselect         (currctrl_sys_register_ram_s2_chipselect),                                    //                                .chipselect
		.currctrl_register_ram_s2_clken              (currctrl_sys_register_ram_s2_clken),                                         //                                .clken
		.currctrl_register_ram_s2_write              (currctrl_sys_register_ram_s2_write),                                         //                                .write
		.currctrl_register_ram_s2_readdata           (currctrl_sys_register_ram_s2_readdata),                                      //                                .readdata
		.currctrl_register_ram_s2_writedata          (currctrl_sys_register_ram_s2_writedata),                                     //                                .writedata
		.currctrl_register_ram_s2_byteenable         (currctrl_sys_register_ram_s2_byteenable),                                    //                                .byteenable
		.currctrlsys_bridge_acknowledge              (currctrl_sys_bridge_acknowledge),                                            //              currctrlsys_bridge.acknowledge
		.currctrlsys_bridge_irq                      (currctrl_sys_bridge_irq),                                                    //                                .irq
		.currctrlsys_bridge_address                  (currctrl_sys_bridge_address),                                                //                                .address
		.currctrlsys_bridge_bus_enable               (currctrl_sys_bridge_bus_enable),                                             //                                .bus_enable
		.currctrlsys_bridge_byte_enable              (currctrl_sys_bridge_byte_enable),                                            //                                .byte_enable
		.currctrlsys_bridge_rw                       (currctrl_sys_bridge_rw),                                                     //                                .rw
		.currctrlsys_bridge_write_data               (currctrl_sys_bridge_write_data),                                             //                                .write_data
		.currctrlsys_bridge_read_data                (currctrl_sys_bridge_read_data),                                              //                                .read_data
		.currctrlsys_bridge_avalon_slave_address     (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_address),     // currctrlsys_bridge_avalon_slave.address
		.currctrlsys_bridge_avalon_slave_byteenable  (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_byteenable),  //                                .byteenable
		.currctrlsys_bridge_avalon_slave_chipselect  (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_chipselect),  //                                .chipselect
		.currctrlsys_bridge_avalon_slave_read        (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_read),        //                                .read
		.currctrlsys_bridge_avalon_slave_write       (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_write),       //                                .write
		.currctrlsys_bridge_avalon_slave_writedata   (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_writedata),   //                                .writedata
		.currctrlsys_bridge_avalon_slave_readdata    (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_readdata),    //                                .readdata
		.currctrlsys_bridge_avalon_slave_waitrequest (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_waitrequest), //                                .waitrequest
		.currctrlsys_bridge_interrupt_irq            (irq_synchronizer_001_receiver_irq),                                          //    currctrlsys_bridge_interrupt.irq
		.reset_currctrl_sys_fifo_reset_n             (reset_currctrl_fifo_reset_n),                                                //         reset_currctrl_sys_fifo.reset_n
		.reset_currctrl_sys_ram_reset_n              (reset_currctrl_ram_reset_n),                                                 //          reset_currctrl_sys_ram.reset_n
		.reset_pheripal_reset_n                      (reset_reset_n)                                                               //                  reset_pheripal.reset_n
	);

	Mk8_InlineController_CPU_Data_Memory data_memory (
		.clk        (altpll_sys_c0_clk),                           //   clk1.clk
		.address    (mm_interconnect_0_data_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_data_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_data_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_data_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_data_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_data_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_data_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze     (1'b0)                                         // (terminated)
	);

	Mk8_InlineController_CPU_Parameter_SYS parameter_sys (
		.clk_ext_ram_clk                                (clk_parameter_ram_clk_clk),                                                //                        clk_ext_ram.clk
		.cpu_clk_clk                                    (altpll_sys_c0_clk),                                                        //                            cpu_clk.clk
		.cpu_reset_reset_n                              (reset_reset_n),                                                            //                          cpu_reset.reset_n
		.crc_init_bridge_avalon_slave_address           (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_address),     //       crc_init_bridge_avalon_slave.address
		.crc_init_bridge_avalon_slave_byteenable        (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_byteenable),  //                                   .byteenable
		.crc_init_bridge_avalon_slave_chipselect        (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_chipselect),  //                                   .chipselect
		.crc_init_bridge_avalon_slave_read              (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_read),        //                                   .read
		.crc_init_bridge_avalon_slave_write             (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_write),       //                                   .write
		.crc_init_bridge_avalon_slave_writedata         (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_writedata),   //                                   .writedata
		.crc_init_bridge_avalon_slave_readdata          (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_readdata),    //                                   .readdata
		.crc_init_bridge_avalon_slave_waitrequest       (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_waitrequest), //                                   .waitrequest
		.crc_init_bridge_external_interface_acknowledge (parameter_sys_crc_init_bridge_acknowledge),                                // crc_init_bridge_external_interface.acknowledge
		.crc_init_bridge_external_interface_irq         (parameter_sys_crc_init_bridge_irq),                                        //                                   .irq
		.crc_init_bridge_external_interface_address     (parameter_sys_crc_init_bridge_address),                                    //                                   .address
		.crc_init_bridge_external_interface_bus_enable  (parameter_sys_crc_init_bridge_bus_enable),                                 //                                   .bus_enable
		.crc_init_bridge_external_interface_byte_enable (parameter_sys_crc_init_bridge_byte_enable),                                //                                   .byte_enable
		.crc_init_bridge_external_interface_rw          (parameter_sys_crc_init_bridge_rw),                                         //                                   .rw
		.crc_init_bridge_external_interface_write_data  (parameter_sys_crc_init_bridge_write_data),                                 //                                   .write_data
		.crc_init_bridge_external_interface_read_data   (parameter_sys_crc_init_bridge_read_data),                                  //                                   .read_data
		.crc_init_bridge_interrupt_irq                  (irq_synchronizer_receiver_irq),                                            //          crc_init_bridge_interrupt.irq
		.parameter_gpio_external_in_port                (parameter_sys_parameter_gpio_in_port),                                     //            parameter_gpio_external.in_port
		.parameter_gpio_external_out_port               (parameter_sys_parameter_gpio_out_port),                                    //                                   .out_port
		.parameter_gpio_s1_address                      (mm_interconnect_1_parameter_sys_parameter_gpio_s1_address),                //                  parameter_gpio_s1.address
		.parameter_gpio_s1_write_n                      (~mm_interconnect_1_parameter_sys_parameter_gpio_s1_write),                 //                                   .write_n
		.parameter_gpio_s1_writedata                    (mm_interconnect_1_parameter_sys_parameter_gpio_s1_writedata),              //                                   .writedata
		.parameter_gpio_s1_chipselect                   (mm_interconnect_1_parameter_sys_parameter_gpio_s1_chipselect),             //                                   .chipselect
		.parameter_gpio_s1_readdata                     (mm_interconnect_1_parameter_sys_parameter_gpio_s1_readdata),               //                                   .readdata
		.parameter_loop_gpio_irq_irq                    (irq_synchronizer_002_receiver_irq),                                        //            parameter_loop_gpio_irq.irq
		.parameter_rx_ram_s1_address                    (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_address),              //                parameter_rx_ram_s1.address
		.parameter_rx_ram_s1_clken                      (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_clken),                //                                   .clken
		.parameter_rx_ram_s1_chipselect                 (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_chipselect),           //                                   .chipselect
		.parameter_rx_ram_s1_write                      (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_write),                //                                   .write
		.parameter_rx_ram_s1_readdata                   (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_readdata),             //                                   .readdata
		.parameter_rx_ram_s1_writedata                  (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_writedata),            //                                   .writedata
		.parameter_rx_ram_s1_byteenable                 (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_byteenable),           //                                   .byteenable
		.parameter_rx_ram_s2_address                    (parameter_sys_parameter_rx_ram_s2_address),                                //                parameter_rx_ram_s2.address
		.parameter_rx_ram_s2_chipselect                 (parameter_sys_parameter_rx_ram_s2_chipselect),                             //                                   .chipselect
		.parameter_rx_ram_s2_clken                      (parameter_sys_parameter_rx_ram_s2_clken),                                  //                                   .clken
		.parameter_rx_ram_s2_write                      (parameter_sys_parameter_rx_ram_s2_write),                                  //                                   .write
		.parameter_rx_ram_s2_readdata                   (parameter_sys_parameter_rx_ram_s2_readdata),                               //                                   .readdata
		.parameter_rx_ram_s2_writedata                  (parameter_sys_parameter_rx_ram_s2_writedata),                              //                                   .writedata
		.parameter_rx_ram_s2_byteenable                 (parameter_sys_parameter_rx_ram_s2_byteenable),                             //                                   .byteenable
		.parameter_tx_ram_s1_address                    (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_address),              //                parameter_tx_ram_s1.address
		.parameter_tx_ram_s1_clken                      (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_clken),                //                                   .clken
		.parameter_tx_ram_s1_chipselect                 (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_chipselect),           //                                   .chipselect
		.parameter_tx_ram_s1_write                      (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_write),                //                                   .write
		.parameter_tx_ram_s1_readdata                   (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_readdata),             //                                   .readdata
		.parameter_tx_ram_s1_writedata                  (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_writedata),            //                                   .writedata
		.parameter_tx_ram_s1_byteenable                 (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_byteenable),           //                                   .byteenable
		.parameter_tx_ram_s2_address                    (parameter_sys_parameter_tx_ram_s2_address),                                //                parameter_tx_ram_s2.address
		.parameter_tx_ram_s2_chipselect                 (parameter_sys_parameter_tx_ram_s2_chipselect),                             //                                   .chipselect
		.parameter_tx_ram_s2_clken                      (parameter_sys_parameter_tx_ram_s2_clken),                                  //                                   .clken
		.parameter_tx_ram_s2_write                      (parameter_sys_parameter_tx_ram_s2_write),                                  //                                   .write
		.parameter_tx_ram_s2_readdata                   (parameter_sys_parameter_tx_ram_s2_readdata),                               //                                   .readdata
		.parameter_tx_ram_s2_writedata                  (parameter_sys_parameter_tx_ram_s2_writedata),                              //                                   .writedata
		.parameter_tx_ram_s2_byteenable                 (parameter_sys_parameter_tx_ram_s2_byteenable),                             //                                   .byteenable
		.parameterlengthpage_export                     (parameter_sys_parameterlengthpage_export),                                 //                parameterlengthpage.export
		.parameterlengthpage_s1_address                 (mm_interconnect_1_parameter_sys_parameterlengthpage_s1_address),           //             parameterlengthpage_s1.address
		.parameterlengthpage_s1_write_n                 (~mm_interconnect_1_parameter_sys_parameterlengthpage_s1_write),            //                                   .write_n
		.parameterlengthpage_s1_writedata               (mm_interconnect_1_parameter_sys_parameterlengthpage_s1_writedata),         //                                   .writedata
		.parameterlengthpage_s1_chipselect              (mm_interconnect_1_parameter_sys_parameterlengthpage_s1_chipselect),        //                                   .chipselect
		.parameterlengthpage_s1_readdata                (mm_interconnect_1_parameter_sys_parameterlengthpage_s1_readdata),          //                                   .readdata
		.pheriphal_clk_clk                              (clk_clk),                                                                  //                      pheriphal_clk.clk
		.pheriphal_reset_reset_n                        (reset_reset_n),                                                            //                    pheriphal_reset.reset_n
		.reset_ext_ram_reset_n                          (reset_parameter_ram_clk_reset_n)                                           //                      reset_ext_ram.reset_n
	);

	Mk8_InlineController_CPU_Pheriphals pheriphals (
		.led_gpio_external_connection_in_port  (pheriphals_led_gpio_external_connection_in_port),     // led_gpio_external_connection.in_port
		.led_gpio_external_connection_out_port (pheriphals_led_gpio_external_connection_out_port),    //                             .out_port
		.led_gpio_s1_address                   (mm_interconnect_1_pheriphals_led_gpio_s1_address),    //                  led_gpio_s1.address
		.led_gpio_s1_write_n                   (~mm_interconnect_1_pheriphals_led_gpio_s1_write),     //                             .write_n
		.led_gpio_s1_writedata                 (mm_interconnect_1_pheriphals_led_gpio_s1_writedata),  //                             .writedata
		.led_gpio_s1_chipselect                (mm_interconnect_1_pheriphals_led_gpio_s1_chipselect), //                             .chipselect
		.led_gpio_s1_readdata                  (mm_interconnect_1_pheriphals_led_gpio_s1_readdata),   //                             .readdata
		.pheriphal_clk_clk                     (clk_clk),                                             //                pheriphal_clk.clk
		.pheriphal_reset_reset_n               (reset_reset_n),                                       //              pheriphal_reset.reset_n
		.tp_gpio_external_connection_export    (pheriphals_tp_gpio_external_connection_export),       //  tp_gpio_external_connection.export
		.tp_gpio_s1_address                    (mm_interconnect_1_pheriphals_tp_gpio_s1_address),     //                   tp_gpio_s1.address
		.tp_gpio_s1_write_n                    (~mm_interconnect_1_pheriphals_tp_gpio_s1_write),      //                             .write_n
		.tp_gpio_s1_writedata                  (mm_interconnect_1_pheriphals_tp_gpio_s1_writedata),   //                             .writedata
		.tp_gpio_s1_chipselect                 (mm_interconnect_1_pheriphals_tp_gpio_s1_chipselect),  //                             .chipselect
		.tp_gpio_s1_readdata                   (mm_interconnect_1_pheriphals_tp_gpio_s1_readdata)     //                             .readdata
	);

	Mk8_InlineController_CPU_Program_Memory program_memory (
		.clk        (altpll_sys_c0_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_program_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_program_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_program_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_program_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_program_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_program_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_program_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	Mk8_InlineController_CPU_TimerSYS timersys (
		.timer_0_irq_irq       (irq_synchronizer_003_receiver_irq),                // timer_0_irq.irq
		.timer_0_s1_address    (mm_interconnect_1_timersys_timer_0_s1_address),    //  timer_0_s1.address
		.timer_0_s1_writedata  (mm_interconnect_1_timersys_timer_0_s1_writedata),  //            .writedata
		.timer_0_s1_readdata   (mm_interconnect_1_timersys_timer_0_s1_readdata),   //            .readdata
		.timer_0_s1_chipselect (mm_interconnect_1_timersys_timer_0_s1_chipselect), //            .chipselect
		.timer_0_s1_write_n    (~mm_interconnect_1_timersys_timer_0_s1_write),     //            .write_n
		.timer_1_irq_irq       (irq_synchronizer_004_receiver_irq),                // timer_1_irq.irq
		.timer_1_s1_address    (mm_interconnect_1_timersys_timer_1_s1_address),    //  timer_1_s1.address
		.timer_1_s1_writedata  (mm_interconnect_1_timersys_timer_1_s1_writedata),  //            .writedata
		.timer_1_s1_readdata   (mm_interconnect_1_timersys_timer_1_s1_readdata),   //            .readdata
		.timer_1_s1_chipselect (mm_interconnect_1_timersys_timer_1_s1_chipselect), //            .chipselect
		.timer_1_s1_write_n    (~mm_interconnect_1_timersys_timer_1_s1_write),     //            .write_n
		.timer_2_irq_irq       (irq_synchronizer_005_receiver_irq),                // timer_2_irq.irq
		.timer_2_s1_address    (mm_interconnect_1_timersys_timer_2_s1_address),    //  timer_2_s1.address
		.timer_2_s1_writedata  (mm_interconnect_1_timersys_timer_2_s1_writedata),  //            .writedata
		.timer_2_s1_readdata   (mm_interconnect_1_timersys_timer_2_s1_readdata),   //            .readdata
		.timer_2_s1_chipselect (mm_interconnect_1_timersys_timer_2_s1_chipselect), //            .chipselect
		.timer_2_s1_write_n    (~mm_interconnect_1_timersys_timer_2_s1_write),     //            .write_n
		.timer_clk_clk         (clk_clk),                                          //   timer_clk.clk
		.timer_reset_reset_n   (reset_reset_n)                                     // timer_reset.reset_n
	);

	Mk8_InlineController_CPU_USB_Data_SYS usb_data_sys (
		.clk_usb_ext_clk_clk        (clk_usb_ext_clk_clk),                                     //   clk_usb_ext_clk.clk
		.cpu_clk_clk                (altpll_sys_c0_clk),                                       //           cpu_clk.clk
		.cpu_reset_reset_n          (reset_reset_n),                                           //         cpu_reset.reset_n
		.pheriphal_clk_clk          (clk_clk),                                                 //     pheriphal_clk.clk
		.pheriphal_reset_reset_n    (reset_reset_n),                                           //   pheriphal_reset.reset_n
		.reset_usb_ext_clk_reset_n  (reset_usb_ext_clk_reset_n),                               // reset_usb_ext_clk.reset_n
		.usb_data_gpio_in_port      (usb_data_sys_usb_data_gpio_in_port),                      //     usb_data_gpio.in_port
		.usb_data_gpio_out_port     (usb_data_sys_usb_data_gpio_out_port),                     //                  .out_port
		.usb_data_gpio_irq_irq      (irq_synchronizer_006_receiver_irq),                       // usb_data_gpio_irq.irq
		.usb_data_ram_s2_address    (usb_data_sys_usb_data_ram_s2_address),                    //   usb_data_ram_s2.address
		.usb_data_ram_s2_chipselect (usb_data_sys_usb_data_ram_s2_chipselect),                 //                  .chipselect
		.usb_data_ram_s2_clken      (usb_data_sys_usb_data_ram_s2_clken),                      //                  .clken
		.usb_data_ram_s2_write      (usb_data_sys_usb_data_ram_s2_write),                      //                  .write
		.usb_data_ram_s2_readdata   (usb_data_sys_usb_data_ram_s2_readdata),                   //                  .readdata
		.usb_data_ram_s2_writedata  (usb_data_sys_usb_data_ram_s2_writedata),                  //                  .writedata
		.usb_data_ram_s2_byteenable (usb_data_sys_usb_data_ram_s2_byteenable),                 //                  .byteenable
		.usb_gpio_s1_address        (mm_interconnect_1_usb_data_sys_usb_gpio_s1_address),      //       usb_gpio_s1.address
		.usb_gpio_s1_write_n        (~mm_interconnect_1_usb_data_sys_usb_gpio_s1_write),       //                  .write_n
		.usb_gpio_s1_writedata      (mm_interconnect_1_usb_data_sys_usb_gpio_s1_writedata),    //                  .writedata
		.usb_gpio_s1_chipselect     (mm_interconnect_1_usb_data_sys_usb_gpio_s1_chipselect),   //                  .chipselect
		.usb_gpio_s1_readdata       (mm_interconnect_1_usb_data_sys_usb_gpio_s1_readdata),     //                  .readdata
		.usb_rx_ram_s1_address      (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_address),    //     usb_rx_ram_s1.address
		.usb_rx_ram_s1_clken        (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_clken),      //                  .clken
		.usb_rx_ram_s1_chipselect   (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_chipselect), //                  .chipselect
		.usb_rx_ram_s1_write        (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_write),      //                  .write
		.usb_rx_ram_s1_readdata     (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_readdata),   //                  .readdata
		.usb_rx_ram_s1_writedata    (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_writedata),  //                  .writedata
		.usb_rx_ram_s1_byteenable   (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_byteenable)  //                  .byteenable
	);

	Mk8_InlineController_CPU_altpll_sys altpll_sys (
		.clk                (clk_clk),                                          //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),               // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_sys_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_sys_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_sys_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_sys_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_sys_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_sys_c0_clk),                                //                    c0.clk
		.c1                 (clk_10m_clk),                                      //                    c1.clk
		.locked             (altpll_sys_locked_conduit_export),                 //        locked_conduit.export
		.scandone           (),                                                 //           (terminated)
		.scandataout        (),                                                 //           (terminated)
		.c2                 (),                                                 //           (terminated)
		.c3                 (),                                                 //           (terminated)
		.c4                 (),                                                 //           (terminated)
		.areset             (1'b0),                                             //           (terminated)
		.phasedone          (),                                                 //           (terminated)
		.phasecounterselect (3'b000),                                           //           (terminated)
		.phaseupdown        (1'b0),                                             //           (terminated)
		.phasestep          (1'b0),                                             //           (terminated)
		.scanclk            (1'b0),                                             //           (terminated)
		.scanclkena         (1'b0),                                             //           (terminated)
		.scandata           (1'b0),                                             //           (terminated)
		.configupdate       (1'b0)                                              //           (terminated)
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (11),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_1 (
		.m0_clk           (clk_clk),                                                       //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                            // m0_reset.reset
		.s0_clk           (altpll_sys_c0_clk),                                             //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                                // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_1_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_1_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_1_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_1_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_1_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_1_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_1_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_1_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_1_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_1_m0_debugaccess)                      //         .debugaccess
	);

	Mk8_InlineController_CPU_msgdma_0 msgdma_0 (
		.mm_read_address              (msgdma_0_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (msgdma_0_mm_read_read),                                   //                 .read
		.mm_read_byteenable           (msgdma_0_mm_read_byteenable),                             //                 .byteenable
		.mm_read_readdata             (msgdma_0_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (msgdma_0_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (msgdma_0_mm_read_readdatavalid),                          //                 .readdatavalid
		.mm_write_address             (msgdma_0_mm_write_address),                               //         mm_write.address
		.mm_write_write               (msgdma_0_mm_write_write),                                 //                 .write
		.mm_write_byteenable          (msgdma_0_mm_write_byteenable),                            //                 .byteenable
		.mm_write_writedata           (msgdma_0_mm_write_writedata),                             //                 .writedata
		.mm_write_waitrequest         (msgdma_0_mm_write_waitrequest),                           //                 .waitrequest
		.clock_clk                    (altpll_sys_c0_clk),                                       //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                         //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_msgdma_0_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_msgdma_0_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_msgdma_0_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_msgdma_0_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_msgdma_0_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_msgdma_0_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_msgdma_0_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_msgdma_0_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_msgdma_0_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_msgdma_0_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_receiver1_irq)                                 //          csr_irq.irq
	);

	Mk8_InlineController_CPU_nios2_gen2 nios2_gen2 (
		.clk                                 (altpll_sys_c0_clk),                                        //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.eic_port_valid                      (vic_0_interrupt_controller_out_valid),                     //   interrupt_controller_in.valid
		.eic_port_data                       (vic_0_interrupt_controller_out_data),                      //                          .data
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (nios2_gen2_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (nios2_gen2_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (nios2_gen2_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (nios2_gen2_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (nios2_gen2_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (nios2_gen2_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (nios2_gen2_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (nios2_gen2_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (nios2_gen2_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (nios2_gen2_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (nios2_gen2_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (nios2_gen2_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (nios2_gen2_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (nios2_gen2_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (nios2_gen2_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (nios2_gen2_custom_instruction_master_multi_writerc),       //                          .multi_writerc
		.E_ci_combo_result                   (nios2_gen2_custom_instruction_master_result),              //                          .result
		.E_ci_combo_a                        (nios2_gen2_custom_instruction_master_a),                   //                          .a
		.E_ci_combo_b                        (nios2_gen2_custom_instruction_master_b),                   //                          .b
		.E_ci_combo_c                        (nios2_gen2_custom_instruction_master_c),                   //                          .c
		.E_ci_combo_dataa                    (nios2_gen2_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_combo_datab                    (nios2_gen2_custom_instruction_master_datab),               //                          .datab
		.E_ci_combo_estatus                  (nios2_gen2_custom_instruction_master_estatus),             //                          .estatus
		.E_ci_combo_ipending                 (nios2_gen2_custom_instruction_master_ipending),            //                          .ipending
		.E_ci_combo_n                        (nios2_gen2_custom_instruction_master_n),                   //                          .n
		.E_ci_combo_readra                   (nios2_gen2_custom_instruction_master_readra),              //                          .readra
		.E_ci_combo_readrb                   (nios2_gen2_custom_instruction_master_readrb),              //                          .readrb
		.E_ci_combo_writerc                  (nios2_gen2_custom_instruction_master_writerc)              //                          .writerc
	);

	Mk8_InlineController_CPU_nios_custom_instr_floating_point_2_0 #(
		.arithmetic_present (1),
		.root_present       (0),
		.conversion_present (1),
		.comparison_present (1)
	) nios_custom_instr_floating_point_2_0 (
		.s1_dataa     (nios2_gen2_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (nios2_gen2_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (nios2_gen2_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (nios2_gen2_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	Mk8_InlineController_CPU_vic_0 vic_0 (
		.clk_clk                        (altpll_sys_c0_clk),                            //                      clk.clk
		.reset_reset                    (rst_controller_reset_out_reset),               //                    reset.reset
		.irq_input_irq                  (vic_0_irq_input_irq),                          //                irq_input.irq
		.csr_access_read                (mm_interconnect_0_vic_0_csr_access_read),      //               csr_access.read
		.csr_access_write               (mm_interconnect_0_vic_0_csr_access_write),     //                         .write
		.csr_access_address             (mm_interconnect_0_vic_0_csr_access_address),   //                         .address
		.csr_access_writedata           (mm_interconnect_0_vic_0_csr_access_writedata), //                         .writedata
		.csr_access_readdata            (mm_interconnect_0_vic_0_csr_access_readdata),  //                         .readdata
		.interrupt_controller_out_valid (vic_0_interrupt_controller_out_valid),         // interrupt_controller_out.valid
		.interrupt_controller_out_data  (vic_0_interrupt_controller_out_data)           //                         .data
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_gen2_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_gen2_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios2_gen2_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios2_gen2_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios2_gen2_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios2_gen2_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios2_gen2_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios2_gen2_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios2_gen2_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios2_gen2_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios2_gen2_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (nios2_gen2_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (nios2_gen2_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (nios2_gen2_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_gen2_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_gen2_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_gen2_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_gen2_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_gen2_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_gen2_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_gen2_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_gen2_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_gen2_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_gen2_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_gen2_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_gen2_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_gen2_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_gen2_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_gen2_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_dataa      (nios2_gen2_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (nios2_gen2_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (nios2_gen2_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (nios2_gen2_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (nios2_gen2_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (nios2_gen2_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (nios2_gen2_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (nios2_gen2_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (nios2_gen2_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (nios2_gen2_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (nios2_gen2_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (nios2_gen2_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (nios2_gen2_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_gen2_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_gen2_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_gen2_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_gen2_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_gen2_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_gen2_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_gen2_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_gen2_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_gen2_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_gen2_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_gen2_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_gen2_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_gen2_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_gen2_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_gen2_custom_instruction_master_translator_multi_ci_master_c)          //                .c
	);

	Mk8_InlineController_CPU_nios2_gen2_custom_instruction_master_comb_xconnect nios2_gen2_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nios2_gen2_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nios2_gen2_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nios2_gen2_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nios2_gen2_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nios2_gen2_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nios2_gen2_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nios2_gen2_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nios2_gen2_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nios2_gen2_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nios2_gen2_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nios2_gen2_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nios2_gen2_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) nios2_gen2_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_gen2_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nios2_gen2_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_gen2_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_gen2_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_gen2_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                             // (terminated)
		.ci_master_readrb    (),                                                                             // (terminated)
		.ci_master_writerc   (),                                                                             // (terminated)
		.ci_master_a         (),                                                                             // (terminated)
		.ci_master_b         (),                                                                             // (terminated)
		.ci_master_c         (),                                                                             // (terminated)
		.ci_master_ipending  (),                                                                             // (terminated)
		.ci_master_estatus   (),                                                                             // (terminated)
		.ci_master_clk       (),                                                                             // (terminated)
		.ci_master_clken     (),                                                                             // (terminated)
		.ci_master_reset_req (),                                                                             // (terminated)
		.ci_master_reset     (),                                                                             // (terminated)
		.ci_master_start     (),                                                                             // (terminated)
		.ci_master_done      (1'b0),                                                                         // (terminated)
		.ci_slave_clk        (1'b0),                                                                         // (terminated)
		.ci_slave_clken      (1'b0),                                                                         // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                         // (terminated)
		.ci_slave_reset      (1'b0),                                                                         // (terminated)
		.ci_slave_start      (1'b0),                                                                         // (terminated)
		.ci_slave_done       ()                                                                              // (terminated)
	);

	Mk8_InlineController_CPU_nios2_gen2_custom_instruction_master_multi_xconnect nios2_gen2_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_gen2_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_gen2_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_gen2_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_gen2_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_gen2_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_gen2_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_gen2_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_gen2_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_gen2_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_gen2_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                          //           .ipending
		.ci_slave_estatus     (),                                                                          //           .estatus
		.ci_slave_clk         (nios2_gen2_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_gen2_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_gen2_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_gen2_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_gen2_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_gen2_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) nios2_gen2_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (nios2_gen2_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (nios2_gen2_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                                 // (terminated)
		.ci_master_readrb    (),                                                                                 // (terminated)
		.ci_master_writerc   (),                                                                                 // (terminated)
		.ci_master_a         (),                                                                                 // (terminated)
		.ci_master_b         (),                                                                                 // (terminated)
		.ci_master_c         (),                                                                                 // (terminated)
		.ci_master_ipending  (),                                                                                 // (terminated)
		.ci_master_estatus   ()                                                                                  // (terminated)
	);

	Mk8_InlineController_CPU_mm_interconnect_0 mm_interconnect_0 (
		.altpll_sys_c0_clk                                            (altpll_sys_c0_clk),                                              //                                          altpll_sys_c0.clk
		.clk_50_clk_clk                                               (clk_clk),                                                        //                                             clk_50_clk.clk
		.altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                             // altpll_sys_inclk_interface_reset_reset_bridge_in_reset.reset
		.msgdma_0_reset_n_reset_bridge_in_reset_reset                 (rst_controller_reset_out_reset),                                 //                 msgdma_0_reset_n_reset_bridge_in_reset.reset
		.nios2_gen2_reset_reset_bridge_in_reset_reset                 (rst_controller_002_reset_out_reset),                             //                 nios2_gen2_reset_reset_bridge_in_reset.reset
		.Parameter_SYS_cpu_reset_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                                 //          Parameter_SYS_cpu_reset_reset_bridge_in_reset.reset
		.msgdma_0_mm_read_address                                     (msgdma_0_mm_read_address),                                       //                                       msgdma_0_mm_read.address
		.msgdma_0_mm_read_waitrequest                                 (msgdma_0_mm_read_waitrequest),                                   //                                                       .waitrequest
		.msgdma_0_mm_read_byteenable                                  (msgdma_0_mm_read_byteenable),                                    //                                                       .byteenable
		.msgdma_0_mm_read_read                                        (msgdma_0_mm_read_read),                                          //                                                       .read
		.msgdma_0_mm_read_readdata                                    (msgdma_0_mm_read_readdata),                                      //                                                       .readdata
		.msgdma_0_mm_read_readdatavalid                               (msgdma_0_mm_read_readdatavalid),                                 //                                                       .readdatavalid
		.msgdma_0_mm_write_address                                    (msgdma_0_mm_write_address),                                      //                                      msgdma_0_mm_write.address
		.msgdma_0_mm_write_waitrequest                                (msgdma_0_mm_write_waitrequest),                                  //                                                       .waitrequest
		.msgdma_0_mm_write_byteenable                                 (msgdma_0_mm_write_byteenable),                                   //                                                       .byteenable
		.msgdma_0_mm_write_write                                      (msgdma_0_mm_write_write),                                        //                                                       .write
		.msgdma_0_mm_write_writedata                                  (msgdma_0_mm_write_writedata),                                    //                                                       .writedata
		.nios2_gen2_data_master_address                               (nios2_gen2_data_master_address),                                 //                                 nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                           (nios2_gen2_data_master_waitrequest),                             //                                                       .waitrequest
		.nios2_gen2_data_master_byteenable                            (nios2_gen2_data_master_byteenable),                              //                                                       .byteenable
		.nios2_gen2_data_master_read                                  (nios2_gen2_data_master_read),                                    //                                                       .read
		.nios2_gen2_data_master_readdata                              (nios2_gen2_data_master_readdata),                                //                                                       .readdata
		.nios2_gen2_data_master_write                                 (nios2_gen2_data_master_write),                                   //                                                       .write
		.nios2_gen2_data_master_writedata                             (nios2_gen2_data_master_writedata),                               //                                                       .writedata
		.nios2_gen2_data_master_debugaccess                           (nios2_gen2_data_master_debugaccess),                             //                                                       .debugaccess
		.nios2_gen2_instruction_master_address                        (nios2_gen2_instruction_master_address),                          //                          nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest                    (nios2_gen2_instruction_master_waitrequest),                      //                                                       .waitrequest
		.nios2_gen2_instruction_master_read                           (nios2_gen2_instruction_master_read),                             //                                                       .read
		.nios2_gen2_instruction_master_readdata                       (nios2_gen2_instruction_master_readdata),                         //                                                       .readdata
		.nios2_gen2_instruction_master_readdatavalid                  (nios2_gen2_instruction_master_readdatavalid),                    //                                                       .readdatavalid
		.altpll_sys_pll_slave_address                                 (mm_interconnect_0_altpll_sys_pll_slave_address),                 //                                   altpll_sys_pll_slave.address
		.altpll_sys_pll_slave_write                                   (mm_interconnect_0_altpll_sys_pll_slave_write),                   //                                                       .write
		.altpll_sys_pll_slave_read                                    (mm_interconnect_0_altpll_sys_pll_slave_read),                    //                                                       .read
		.altpll_sys_pll_slave_readdata                                (mm_interconnect_0_altpll_sys_pll_slave_readdata),                //                                                       .readdata
		.altpll_sys_pll_slave_writedata                               (mm_interconnect_0_altpll_sys_pll_slave_writedata),               //                                                       .writedata
		.Data_Memory_s1_address                                       (mm_interconnect_0_data_memory_s1_address),                       //                                         Data_Memory_s1.address
		.Data_Memory_s1_write                                         (mm_interconnect_0_data_memory_s1_write),                         //                                                       .write
		.Data_Memory_s1_readdata                                      (mm_interconnect_0_data_memory_s1_readdata),                      //                                                       .readdata
		.Data_Memory_s1_writedata                                     (mm_interconnect_0_data_memory_s1_writedata),                     //                                                       .writedata
		.Data_Memory_s1_byteenable                                    (mm_interconnect_0_data_memory_s1_byteenable),                    //                                                       .byteenable
		.Data_Memory_s1_chipselect                                    (mm_interconnect_0_data_memory_s1_chipselect),                    //                                                       .chipselect
		.Data_Memory_s1_clken                                         (mm_interconnect_0_data_memory_s1_clken),                         //                                                       .clken
		.mm_clock_crossing_bridge_1_s0_address                        (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_address),        //                          mm_clock_crossing_bridge_1_s0.address
		.mm_clock_crossing_bridge_1_s0_write                          (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_write),          //                                                       .write
		.mm_clock_crossing_bridge_1_s0_read                           (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_read),           //                                                       .read
		.mm_clock_crossing_bridge_1_s0_readdata                       (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdata),       //                                                       .readdata
		.mm_clock_crossing_bridge_1_s0_writedata                      (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_writedata),      //                                                       .writedata
		.mm_clock_crossing_bridge_1_s0_burstcount                     (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_burstcount),     //                                                       .burstcount
		.mm_clock_crossing_bridge_1_s0_byteenable                     (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_byteenable),     //                                                       .byteenable
		.mm_clock_crossing_bridge_1_s0_readdatavalid                  (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdatavalid),  //                                                       .readdatavalid
		.mm_clock_crossing_bridge_1_s0_waitrequest                    (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_waitrequest),    //                                                       .waitrequest
		.mm_clock_crossing_bridge_1_s0_debugaccess                    (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_debugaccess),    //                                                       .debugaccess
		.msgdma_0_csr_address                                         (mm_interconnect_0_msgdma_0_csr_address),                         //                                           msgdma_0_csr.address
		.msgdma_0_csr_write                                           (mm_interconnect_0_msgdma_0_csr_write),                           //                                                       .write
		.msgdma_0_csr_read                                            (mm_interconnect_0_msgdma_0_csr_read),                            //                                                       .read
		.msgdma_0_csr_readdata                                        (mm_interconnect_0_msgdma_0_csr_readdata),                        //                                                       .readdata
		.msgdma_0_csr_writedata                                       (mm_interconnect_0_msgdma_0_csr_writedata),                       //                                                       .writedata
		.msgdma_0_csr_byteenable                                      (mm_interconnect_0_msgdma_0_csr_byteenable),                      //                                                       .byteenable
		.msgdma_0_descriptor_slave_write                              (mm_interconnect_0_msgdma_0_descriptor_slave_write),              //                              msgdma_0_descriptor_slave.write
		.msgdma_0_descriptor_slave_writedata                          (mm_interconnect_0_msgdma_0_descriptor_slave_writedata),          //                                                       .writedata
		.msgdma_0_descriptor_slave_byteenable                         (mm_interconnect_0_msgdma_0_descriptor_slave_byteenable),         //                                                       .byteenable
		.msgdma_0_descriptor_slave_waitrequest                        (mm_interconnect_0_msgdma_0_descriptor_slave_waitrequest),        //                                                       .waitrequest
		.nios2_gen2_debug_mem_slave_address                           (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),           //                             nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                             (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),             //                                                       .write
		.nios2_gen2_debug_mem_slave_read                              (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),              //                                                       .read
		.nios2_gen2_debug_mem_slave_readdata                          (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),          //                                                       .readdata
		.nios2_gen2_debug_mem_slave_writedata                         (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),         //                                                       .writedata
		.nios2_gen2_debug_mem_slave_byteenable                        (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),        //                                                       .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest                       (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),       //                                                       .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess                       (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),       //                                                       .debugaccess
		.Parameter_SYS_parameter_rx_ram_s1_address                    (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_address),    //                      Parameter_SYS_parameter_rx_ram_s1.address
		.Parameter_SYS_parameter_rx_ram_s1_write                      (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_write),      //                                                       .write
		.Parameter_SYS_parameter_rx_ram_s1_readdata                   (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_readdata),   //                                                       .readdata
		.Parameter_SYS_parameter_rx_ram_s1_writedata                  (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_writedata),  //                                                       .writedata
		.Parameter_SYS_parameter_rx_ram_s1_byteenable                 (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_byteenable), //                                                       .byteenable
		.Parameter_SYS_parameter_rx_ram_s1_chipselect                 (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_chipselect), //                                                       .chipselect
		.Parameter_SYS_parameter_rx_ram_s1_clken                      (mm_interconnect_0_parameter_sys_parameter_rx_ram_s1_clken),      //                                                       .clken
		.Parameter_SYS_parameter_tx_ram_s1_address                    (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_address),    //                      Parameter_SYS_parameter_tx_ram_s1.address
		.Parameter_SYS_parameter_tx_ram_s1_write                      (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_write),      //                                                       .write
		.Parameter_SYS_parameter_tx_ram_s1_readdata                   (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_readdata),   //                                                       .readdata
		.Parameter_SYS_parameter_tx_ram_s1_writedata                  (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_writedata),  //                                                       .writedata
		.Parameter_SYS_parameter_tx_ram_s1_byteenable                 (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_byteenable), //                                                       .byteenable
		.Parameter_SYS_parameter_tx_ram_s1_chipselect                 (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_chipselect), //                                                       .chipselect
		.Parameter_SYS_parameter_tx_ram_s1_clken                      (mm_interconnect_0_parameter_sys_parameter_tx_ram_s1_clken),      //                                                       .clken
		.Program_Memory_s1_address                                    (mm_interconnect_0_program_memory_s1_address),                    //                                      Program_Memory_s1.address
		.Program_Memory_s1_write                                      (mm_interconnect_0_program_memory_s1_write),                      //                                                       .write
		.Program_Memory_s1_readdata                                   (mm_interconnect_0_program_memory_s1_readdata),                   //                                                       .readdata
		.Program_Memory_s1_writedata                                  (mm_interconnect_0_program_memory_s1_writedata),                  //                                                       .writedata
		.Program_Memory_s1_byteenable                                 (mm_interconnect_0_program_memory_s1_byteenable),                 //                                                       .byteenable
		.Program_Memory_s1_chipselect                                 (mm_interconnect_0_program_memory_s1_chipselect),                 //                                                       .chipselect
		.Program_Memory_s1_clken                                      (mm_interconnect_0_program_memory_s1_clken),                      //                                                       .clken
		.USB_Data_SYS_usb_rx_ram_s1_address                           (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_address),           //                             USB_Data_SYS_usb_rx_ram_s1.address
		.USB_Data_SYS_usb_rx_ram_s1_write                             (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_write),             //                                                       .write
		.USB_Data_SYS_usb_rx_ram_s1_readdata                          (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_readdata),          //                                                       .readdata
		.USB_Data_SYS_usb_rx_ram_s1_writedata                         (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_writedata),         //                                                       .writedata
		.USB_Data_SYS_usb_rx_ram_s1_byteenable                        (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_byteenable),        //                                                       .byteenable
		.USB_Data_SYS_usb_rx_ram_s1_chipselect                        (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_chipselect),        //                                                       .chipselect
		.USB_Data_SYS_usb_rx_ram_s1_clken                             (mm_interconnect_0_usb_data_sys_usb_rx_ram_s1_clken),             //                                                       .clken
		.vic_0_csr_access_address                                     (mm_interconnect_0_vic_0_csr_access_address),                     //                                       vic_0_csr_access.address
		.vic_0_csr_access_write                                       (mm_interconnect_0_vic_0_csr_access_write),                       //                                                       .write
		.vic_0_csr_access_read                                        (mm_interconnect_0_vic_0_csr_access_read),                        //                                                       .read
		.vic_0_csr_access_readdata                                    (mm_interconnect_0_vic_0_csr_access_readdata),                    //                                                       .readdata
		.vic_0_csr_access_writedata                                   (mm_interconnect_0_vic_0_csr_access_writedata)                    //                                                       .writedata
	);

	Mk8_InlineController_CPU_mm_interconnect_1 mm_interconnect_1 (
		.clk_50_clk_clk                                                  (clk_clk),                                                                    //                                                clk_50_clk.clk
		.mm_clock_crossing_bridge_1_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                         // mm_clock_crossing_bridge_1_m0_reset_reset_bridge_in_reset.reset
		.Parameter_SYS_pheriphal_reset_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),                                         //       Parameter_SYS_pheriphal_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_1_m0_address                           (mm_clock_crossing_bridge_1_m0_address),                                      //                             mm_clock_crossing_bridge_1_m0.address
		.mm_clock_crossing_bridge_1_m0_waitrequest                       (mm_clock_crossing_bridge_1_m0_waitrequest),                                  //                                                          .waitrequest
		.mm_clock_crossing_bridge_1_m0_burstcount                        (mm_clock_crossing_bridge_1_m0_burstcount),                                   //                                                          .burstcount
		.mm_clock_crossing_bridge_1_m0_byteenable                        (mm_clock_crossing_bridge_1_m0_byteenable),                                   //                                                          .byteenable
		.mm_clock_crossing_bridge_1_m0_read                              (mm_clock_crossing_bridge_1_m0_read),                                         //                                                          .read
		.mm_clock_crossing_bridge_1_m0_readdata                          (mm_clock_crossing_bridge_1_m0_readdata),                                     //                                                          .readdata
		.mm_clock_crossing_bridge_1_m0_readdatavalid                     (mm_clock_crossing_bridge_1_m0_readdatavalid),                                //                                                          .readdatavalid
		.mm_clock_crossing_bridge_1_m0_write                             (mm_clock_crossing_bridge_1_m0_write),                                        //                                                          .write
		.mm_clock_crossing_bridge_1_m0_writedata                         (mm_clock_crossing_bridge_1_m0_writedata),                                    //                                                          .writedata
		.mm_clock_crossing_bridge_1_m0_debugaccess                       (mm_clock_crossing_bridge_1_m0_debugaccess),                                  //                                                          .debugaccess
		.CurrCTRL_SYS_currctrl_gpio_s1_address                           (mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_address),                    //                             CurrCTRL_SYS_currctrl_gpio_s1.address
		.CurrCTRL_SYS_currctrl_gpio_s1_write                             (mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_write),                      //                                                          .write
		.CurrCTRL_SYS_currctrl_gpio_s1_readdata                          (mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_readdata),                   //                                                          .readdata
		.CurrCTRL_SYS_currctrl_gpio_s1_writedata                         (mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_writedata),                  //                                                          .writedata
		.CurrCTRL_SYS_currctrl_gpio_s1_chipselect                        (mm_interconnect_1_currctrl_sys_currctrl_gpio_s1_chipselect),                 //                                                          .chipselect
		.CurrCTRL_SYS_currctrl_register_ram_s1_address                   (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_address),            //                     CurrCTRL_SYS_currctrl_register_ram_s1.address
		.CurrCTRL_SYS_currctrl_register_ram_s1_write                     (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_write),              //                                                          .write
		.CurrCTRL_SYS_currctrl_register_ram_s1_readdata                  (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_readdata),           //                                                          .readdata
		.CurrCTRL_SYS_currctrl_register_ram_s1_writedata                 (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_writedata),          //                                                          .writedata
		.CurrCTRL_SYS_currctrl_register_ram_s1_byteenable                (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_byteenable),         //                                                          .byteenable
		.CurrCTRL_SYS_currctrl_register_ram_s1_chipselect                (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_chipselect),         //                                                          .chipselect
		.CurrCTRL_SYS_currctrl_register_ram_s1_clken                     (mm_interconnect_1_currctrl_sys_currctrl_register_ram_s1_clken),              //                                                          .clken
		.CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_address            (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_address),     //              CurrCTRL_SYS_currctrlsys_bridge_avalon_slave.address
		.CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_write              (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_write),       //                                                          .write
		.CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_read               (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_read),        //                                                          .read
		.CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_readdata           (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_readdata),    //                                                          .readdata
		.CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_writedata          (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_writedata),   //                                                          .writedata
		.CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_byteenable         (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_byteenable),  //                                                          .byteenable
		.CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_waitrequest        (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_waitrequest), //                                                          .waitrequest
		.CurrCTRL_SYS_currctrlsys_bridge_avalon_slave_chipselect         (mm_interconnect_1_currctrl_sys_currctrlsys_bridge_avalon_slave_chipselect),  //                                                          .chipselect
		.Parameter_SYS_crc_init_bridge_avalon_slave_address              (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_address),       //                Parameter_SYS_crc_init_bridge_avalon_slave.address
		.Parameter_SYS_crc_init_bridge_avalon_slave_write                (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_write),         //                                                          .write
		.Parameter_SYS_crc_init_bridge_avalon_slave_read                 (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_read),          //                                                          .read
		.Parameter_SYS_crc_init_bridge_avalon_slave_readdata             (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_readdata),      //                                                          .readdata
		.Parameter_SYS_crc_init_bridge_avalon_slave_writedata            (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_writedata),     //                                                          .writedata
		.Parameter_SYS_crc_init_bridge_avalon_slave_byteenable           (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_byteenable),    //                                                          .byteenable
		.Parameter_SYS_crc_init_bridge_avalon_slave_waitrequest          (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_waitrequest),   //                                                          .waitrequest
		.Parameter_SYS_crc_init_bridge_avalon_slave_chipselect           (mm_interconnect_1_parameter_sys_crc_init_bridge_avalon_slave_chipselect),    //                                                          .chipselect
		.Parameter_SYS_parameter_gpio_s1_address                         (mm_interconnect_1_parameter_sys_parameter_gpio_s1_address),                  //                           Parameter_SYS_parameter_gpio_s1.address
		.Parameter_SYS_parameter_gpio_s1_write                           (mm_interconnect_1_parameter_sys_parameter_gpio_s1_write),                    //                                                          .write
		.Parameter_SYS_parameter_gpio_s1_readdata                        (mm_interconnect_1_parameter_sys_parameter_gpio_s1_readdata),                 //                                                          .readdata
		.Parameter_SYS_parameter_gpio_s1_writedata                       (mm_interconnect_1_parameter_sys_parameter_gpio_s1_writedata),                //                                                          .writedata
		.Parameter_SYS_parameter_gpio_s1_chipselect                      (mm_interconnect_1_parameter_sys_parameter_gpio_s1_chipselect),               //                                                          .chipselect
		.Parameter_SYS_parameterlengthpage_s1_address                    (mm_interconnect_1_parameter_sys_parameterlengthpage_s1_address),             //                      Parameter_SYS_parameterlengthpage_s1.address
		.Parameter_SYS_parameterlengthpage_s1_write                      (mm_interconnect_1_parameter_sys_parameterlengthpage_s1_write),               //                                                          .write
		.Parameter_SYS_parameterlengthpage_s1_readdata                   (mm_interconnect_1_parameter_sys_parameterlengthpage_s1_readdata),            //                                                          .readdata
		.Parameter_SYS_parameterlengthpage_s1_writedata                  (mm_interconnect_1_parameter_sys_parameterlengthpage_s1_writedata),           //                                                          .writedata
		.Parameter_SYS_parameterlengthpage_s1_chipselect                 (mm_interconnect_1_parameter_sys_parameterlengthpage_s1_chipselect),          //                                                          .chipselect
		.Pheriphals_led_gpio_s1_address                                  (mm_interconnect_1_pheriphals_led_gpio_s1_address),                           //                                    Pheriphals_led_gpio_s1.address
		.Pheriphals_led_gpio_s1_write                                    (mm_interconnect_1_pheriphals_led_gpio_s1_write),                             //                                                          .write
		.Pheriphals_led_gpio_s1_readdata                                 (mm_interconnect_1_pheriphals_led_gpio_s1_readdata),                          //                                                          .readdata
		.Pheriphals_led_gpio_s1_writedata                                (mm_interconnect_1_pheriphals_led_gpio_s1_writedata),                         //                                                          .writedata
		.Pheriphals_led_gpio_s1_chipselect                               (mm_interconnect_1_pheriphals_led_gpio_s1_chipselect),                        //                                                          .chipselect
		.Pheriphals_tp_gpio_s1_address                                   (mm_interconnect_1_pheriphals_tp_gpio_s1_address),                            //                                     Pheriphals_tp_gpio_s1.address
		.Pheriphals_tp_gpio_s1_write                                     (mm_interconnect_1_pheriphals_tp_gpio_s1_write),                              //                                                          .write
		.Pheriphals_tp_gpio_s1_readdata                                  (mm_interconnect_1_pheriphals_tp_gpio_s1_readdata),                           //                                                          .readdata
		.Pheriphals_tp_gpio_s1_writedata                                 (mm_interconnect_1_pheriphals_tp_gpio_s1_writedata),                          //                                                          .writedata
		.Pheriphals_tp_gpio_s1_chipselect                                (mm_interconnect_1_pheriphals_tp_gpio_s1_chipselect),                         //                                                          .chipselect
		.TimerSYS_timer_0_s1_address                                     (mm_interconnect_1_timersys_timer_0_s1_address),                              //                                       TimerSYS_timer_0_s1.address
		.TimerSYS_timer_0_s1_write                                       (mm_interconnect_1_timersys_timer_0_s1_write),                                //                                                          .write
		.TimerSYS_timer_0_s1_readdata                                    (mm_interconnect_1_timersys_timer_0_s1_readdata),                             //                                                          .readdata
		.TimerSYS_timer_0_s1_writedata                                   (mm_interconnect_1_timersys_timer_0_s1_writedata),                            //                                                          .writedata
		.TimerSYS_timer_0_s1_chipselect                                  (mm_interconnect_1_timersys_timer_0_s1_chipselect),                           //                                                          .chipselect
		.TimerSYS_timer_1_s1_address                                     (mm_interconnect_1_timersys_timer_1_s1_address),                              //                                       TimerSYS_timer_1_s1.address
		.TimerSYS_timer_1_s1_write                                       (mm_interconnect_1_timersys_timer_1_s1_write),                                //                                                          .write
		.TimerSYS_timer_1_s1_readdata                                    (mm_interconnect_1_timersys_timer_1_s1_readdata),                             //                                                          .readdata
		.TimerSYS_timer_1_s1_writedata                                   (mm_interconnect_1_timersys_timer_1_s1_writedata),                            //                                                          .writedata
		.TimerSYS_timer_1_s1_chipselect                                  (mm_interconnect_1_timersys_timer_1_s1_chipselect),                           //                                                          .chipselect
		.TimerSYS_timer_2_s1_address                                     (mm_interconnect_1_timersys_timer_2_s1_address),                              //                                       TimerSYS_timer_2_s1.address
		.TimerSYS_timer_2_s1_write                                       (mm_interconnect_1_timersys_timer_2_s1_write),                                //                                                          .write
		.TimerSYS_timer_2_s1_readdata                                    (mm_interconnect_1_timersys_timer_2_s1_readdata),                             //                                                          .readdata
		.TimerSYS_timer_2_s1_writedata                                   (mm_interconnect_1_timersys_timer_2_s1_writedata),                            //                                                          .writedata
		.TimerSYS_timer_2_s1_chipselect                                  (mm_interconnect_1_timersys_timer_2_s1_chipselect),                           //                                                          .chipselect
		.USB_Data_SYS_usb_gpio_s1_address                                (mm_interconnect_1_usb_data_sys_usb_gpio_s1_address),                         //                                  USB_Data_SYS_usb_gpio_s1.address
		.USB_Data_SYS_usb_gpio_s1_write                                  (mm_interconnect_1_usb_data_sys_usb_gpio_s1_write),                           //                                                          .write
		.USB_Data_SYS_usb_gpio_s1_readdata                               (mm_interconnect_1_usb_data_sys_usb_gpio_s1_readdata),                        //                                                          .readdata
		.USB_Data_SYS_usb_gpio_s1_writedata                              (mm_interconnect_1_usb_data_sys_usb_gpio_s1_writedata),                       //                                                          .writedata
		.USB_Data_SYS_usb_gpio_s1_chipselect                             (mm_interconnect_1_usb_data_sys_usb_gpio_s1_chipselect)                       //                                                          .chipselect
	);

	Mk8_InlineController_CPU_irq_mapper irq_mapper (
		.clk           (altpll_sys_c0_clk),              //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.sender_irq    (vic_0_irq_input_irq)             //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_sys_c0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_sys_c0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_sys_c0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_sys_c0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_sys_c0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver5_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_005 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_sys_c0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_005_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver6_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_006 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_sys_c0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_006_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver7_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (altpll_sys_c0_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset),   // reset_in1.reset
		.clk            (altpll_sys_c0_clk),                      //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	assign cpu_clk_clk = clk_clk;

endmodule
