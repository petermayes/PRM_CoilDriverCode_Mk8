// Pararameter_Comms_SYS.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module Pararameter_Comms_SYS (
		input  wire        clk_ext_ram_clk,                                //                        clk_ext_ram.clk
		input  wire        cpu_clk_clk,                                    //                            cpu_clk.clk
		input  wire        cpu_reset_reset_n,                              //                          cpu_reset.reset_n
		input  wire [7:0]  crc_init_bridge_avalon_slave_address,           //       crc_init_bridge_avalon_slave.address
		input  wire        crc_init_bridge_avalon_slave_byteenable,        //                                   .byteenable
		input  wire        crc_init_bridge_avalon_slave_chipselect,        //                                   .chipselect
		input  wire        crc_init_bridge_avalon_slave_read,              //                                   .read
		input  wire        crc_init_bridge_avalon_slave_write,             //                                   .write
		input  wire [7:0]  crc_init_bridge_avalon_slave_writedata,         //                                   .writedata
		output wire [7:0]  crc_init_bridge_avalon_slave_readdata,          //                                   .readdata
		output wire        crc_init_bridge_avalon_slave_waitrequest,       //                                   .waitrequest
		input  wire        crc_init_bridge_external_interface_acknowledge, // crc_init_bridge_external_interface.acknowledge
		input  wire        crc_init_bridge_external_interface_irq,         //                                   .irq
		output wire [7:0]  crc_init_bridge_external_interface_address,     //                                   .address
		output wire        crc_init_bridge_external_interface_bus_enable,  //                                   .bus_enable
		output wire        crc_init_bridge_external_interface_byte_enable, //                                   .byte_enable
		output wire        crc_init_bridge_external_interface_rw,          //                                   .rw
		output wire [7:0]  crc_init_bridge_external_interface_write_data,  //                                   .write_data
		input  wire [7:0]  crc_init_bridge_external_interface_read_data,   //                                   .read_data
		output wire        crc_init_bridge_interrupt_irq,                  //          crc_init_bridge_interrupt.irq
		input  wire        parameter_gpio_external_in_port,                //            parameter_gpio_external.in_port
		output wire        parameter_gpio_external_out_port,               //                                   .out_port
		input  wire [2:0]  parameter_gpio_s1_address,                      //                  parameter_gpio_s1.address
		input  wire        parameter_gpio_s1_write_n,                      //                                   .write_n
		input  wire [31:0] parameter_gpio_s1_writedata,                    //                                   .writedata
		input  wire        parameter_gpio_s1_chipselect,                   //                                   .chipselect
		output wire [31:0] parameter_gpio_s1_readdata,                     //                                   .readdata
		output wire        parameter_loop_gpio_irq_irq,                    //            parameter_loop_gpio_irq.irq
		input  wire [10:0] parameter_rx_ram_s1_address,                    //                parameter_rx_ram_s1.address
		input  wire        parameter_rx_ram_s1_clken,                      //                                   .clken
		input  wire        parameter_rx_ram_s1_chipselect,                 //                                   .chipselect
		input  wire        parameter_rx_ram_s1_write,                      //                                   .write
		output wire [31:0] parameter_rx_ram_s1_readdata,                   //                                   .readdata
		input  wire [31:0] parameter_rx_ram_s1_writedata,                  //                                   .writedata
		input  wire [3:0]  parameter_rx_ram_s1_byteenable,                 //                                   .byteenable
		input  wire [10:0] parameter_rx_ram_s2_address,                    //                parameter_rx_ram_s2.address
		input  wire        parameter_rx_ram_s2_chipselect,                 //                                   .chipselect
		input  wire        parameter_rx_ram_s2_clken,                      //                                   .clken
		input  wire        parameter_rx_ram_s2_write,                      //                                   .write
		output wire [31:0] parameter_rx_ram_s2_readdata,                   //                                   .readdata
		input  wire [31:0] parameter_rx_ram_s2_writedata,                  //                                   .writedata
		input  wire [3:0]  parameter_rx_ram_s2_byteenable,                 //                                   .byteenable
		input  wire [10:0] parameter_tx_ram_s1_address,                    //                parameter_tx_ram_s1.address
		input  wire        parameter_tx_ram_s1_clken,                      //                                   .clken
		input  wire        parameter_tx_ram_s1_chipselect,                 //                                   .chipselect
		input  wire        parameter_tx_ram_s1_write,                      //                                   .write
		output wire [31:0] parameter_tx_ram_s1_readdata,                   //                                   .readdata
		input  wire [31:0] parameter_tx_ram_s1_writedata,                  //                                   .writedata
		input  wire [3:0]  parameter_tx_ram_s1_byteenable,                 //                                   .byteenable
		input  wire [10:0] parameter_tx_ram_s2_address,                    //                parameter_tx_ram_s2.address
		input  wire        parameter_tx_ram_s2_chipselect,                 //                                   .chipselect
		input  wire        parameter_tx_ram_s2_clken,                      //                                   .clken
		input  wire        parameter_tx_ram_s2_write,                      //                                   .write
		output wire [31:0] parameter_tx_ram_s2_readdata,                   //                                   .readdata
		input  wire [31:0] parameter_tx_ram_s2_writedata,                  //                                   .writedata
		input  wire [3:0]  parameter_tx_ram_s2_byteenable,                 //                                   .byteenable
		output wire [15:0] parameterlengthpage_export,                     //                parameterlengthpage.export
		input  wire [1:0]  parameterlengthpage_s1_address,                 //             parameterlengthpage_s1.address
		input  wire        parameterlengthpage_s1_write_n,                 //                                   .write_n
		input  wire [31:0] parameterlengthpage_s1_writedata,               //                                   .writedata
		input  wire        parameterlengthpage_s1_chipselect,              //                                   .chipselect
		output wire [31:0] parameterlengthpage_s1_readdata,                //                                   .readdata
		input  wire        pheriphal_clk_clk,                              //                      pheriphal_clk.clk
		input  wire        pheriphal_reset_reset_n,                        //                    pheriphal_reset.reset_n
		input  wire        reset_ext_ram_reset_n                           //                      reset_ext_ram.reset_n
	);

	wire    rst_controller_reset_out_reset;         // rst_controller:reset_out -> [CRC_Init_Bridge:reset, ParameterLengthPage:reset_n, Parameter_GPIO:reset_n]
	wire    rst_controller_001_reset_out_reset;     // rst_controller_001:reset_out -> [Parameter_RX_RAM:reset, Parameter_TX_RAM:reset]
	wire    rst_controller_001_reset_out_reset_req; // rst_controller_001:reset_req -> [Parameter_RX_RAM:reset_req, Parameter_TX_RAM:reset_req]
	wire    rst_controller_002_reset_out_reset;     // rst_controller_002:reset_out -> [Parameter_RX_RAM:reset2, Parameter_TX_RAM:reset2]
	wire    rst_controller_002_reset_out_reset_req; // rst_controller_002:reset_req -> [Parameter_RX_RAM:reset_req2, Parameter_TX_RAM:reset_req2]

	Pararameter_Comms_SYS_CRC_Init_Bridge crc_init_bridge (
		.clk                (pheriphal_clk_clk),                              //                clk.clk
		.reset              (rst_controller_reset_out_reset),                 //              reset.reset
		.avalon_address     (crc_init_bridge_avalon_slave_address),           //       avalon_slave.address
		.avalon_byteenable  (crc_init_bridge_avalon_slave_byteenable),        //                   .byteenable
		.avalon_chipselect  (crc_init_bridge_avalon_slave_chipselect),        //                   .chipselect
		.avalon_read        (crc_init_bridge_avalon_slave_read),              //                   .read
		.avalon_write       (crc_init_bridge_avalon_slave_write),             //                   .write
		.avalon_writedata   (crc_init_bridge_avalon_slave_writedata),         //                   .writedata
		.avalon_readdata    (crc_init_bridge_avalon_slave_readdata),          //                   .readdata
		.avalon_waitrequest (crc_init_bridge_avalon_slave_waitrequest),       //                   .waitrequest
		.avalon_irq         (crc_init_bridge_interrupt_irq),                  //          interrupt.irq
		.acknowledge        (crc_init_bridge_external_interface_acknowledge), // external_interface.export
		.irq                (crc_init_bridge_external_interface_irq),         //                   .export
		.address            (crc_init_bridge_external_interface_address),     //                   .export
		.bus_enable         (crc_init_bridge_external_interface_bus_enable),  //                   .export
		.byte_enable        (crc_init_bridge_external_interface_byte_enable), //                   .export
		.rw                 (crc_init_bridge_external_interface_rw),          //                   .export
		.write_data         (crc_init_bridge_external_interface_write_data),  //                   .export
		.read_data          (crc_init_bridge_external_interface_read_data)    //                   .export
	);

	Pararameter_Comms_SYS_ParameterLengthPage parameterlengthpage (
		.clk        (pheriphal_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address    (parameterlengthpage_s1_address),    //                  s1.address
		.write_n    (parameterlengthpage_s1_write_n),    //                    .write_n
		.writedata  (parameterlengthpage_s1_writedata),  //                    .writedata
		.chipselect (parameterlengthpage_s1_chipselect), //                    .chipselect
		.readdata   (parameterlengthpage_s1_readdata),   //                    .readdata
		.out_port   (parameterlengthpage_export)         // external_connection.export
	);

	Pararameter_Comms_SYS_Parameter_GPIO parameter_gpio (
		.clk        (pheriphal_clk_clk),                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address    (parameter_gpio_s1_address),        //                  s1.address
		.write_n    (parameter_gpio_s1_write_n),        //                    .write_n
		.writedata  (parameter_gpio_s1_writedata),      //                    .writedata
		.chipselect (parameter_gpio_s1_chipselect),     //                    .chipselect
		.readdata   (parameter_gpio_s1_readdata),       //                    .readdata
		.in_port    (parameter_gpio_external_in_port),  // external_connection.export
		.out_port   (parameter_gpio_external_out_port), //                    .export
		.irq        (parameter_loop_gpio_irq_irq)       //                 irq.irq
	);

	Pararameter_Comms_SYS_Parameter_RX_RAM parameter_rx_ram (
		.clk         (cpu_clk_clk),                            //   clk1.clk
		.address     (parameter_rx_ram_s1_address),            //     s1.address
		.clken       (parameter_rx_ram_s1_clken),              //       .clken
		.chipselect  (parameter_rx_ram_s1_chipselect),         //       .chipselect
		.write       (parameter_rx_ram_s1_write),              //       .write
		.readdata    (parameter_rx_ram_s1_readdata),           //       .readdata
		.writedata   (parameter_rx_ram_s1_writedata),          //       .writedata
		.byteenable  (parameter_rx_ram_s1_byteenable),         //       .byteenable
		.reset       (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req), //       .reset_req
		.address2    (parameter_rx_ram_s2_address),            //     s2.address
		.chipselect2 (parameter_rx_ram_s2_chipselect),         //       .chipselect
		.clken2      (parameter_rx_ram_s2_clken),              //       .clken
		.write2      (parameter_rx_ram_s2_write),              //       .write
		.readdata2   (parameter_rx_ram_s2_readdata),           //       .readdata
		.writedata2  (parameter_rx_ram_s2_writedata),          //       .writedata
		.byteenable2 (parameter_rx_ram_s2_byteenable),         //       .byteenable
		.clk2        (clk_ext_ram_clk),                        //   clk2.clk
		.reset2      (rst_controller_002_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_002_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	Pararameter_Comms_SYS_Parameter_TX_RAM parameter_tx_ram (
		.clk         (cpu_clk_clk),                            //   clk1.clk
		.address     (parameter_tx_ram_s1_address),            //     s1.address
		.clken       (parameter_tx_ram_s1_clken),              //       .clken
		.chipselect  (parameter_tx_ram_s1_chipselect),         //       .chipselect
		.write       (parameter_tx_ram_s1_write),              //       .write
		.readdata    (parameter_tx_ram_s1_readdata),           //       .readdata
		.writedata   (parameter_tx_ram_s1_writedata),          //       .writedata
		.byteenable  (parameter_tx_ram_s1_byteenable),         //       .byteenable
		.reset       (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req), //       .reset_req
		.address2    (parameter_tx_ram_s2_address),            //     s2.address
		.chipselect2 (parameter_tx_ram_s2_chipselect),         //       .chipselect
		.clken2      (parameter_tx_ram_s2_clken),              //       .clken
		.write2      (parameter_tx_ram_s2_write),              //       .write
		.readdata2   (parameter_tx_ram_s2_readdata),           //       .readdata
		.writedata2  (parameter_tx_ram_s2_writedata),          //       .writedata
		.byteenable2 (parameter_tx_ram_s2_byteenable),         //       .byteenable
		.clk2        (clk_ext_ram_clk),                        //   clk2.clk
		.reset2      (rst_controller_002_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_002_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~pheriphal_reset_reset_n),       // reset_in0.reset
		.clk            (pheriphal_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~cpu_reset_reset_n),                     // reset_in0.reset
		.clk            (cpu_clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_ext_ram_reset_n),                 // reset_in0.reset
		.clk            (clk_ext_ram_clk),                        //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
